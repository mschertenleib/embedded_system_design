module biosRom ( input wire        clock,
                 input wire [10:0] address,
                 output reg [31:0] romData);

  always @(negedge clock)
    case (address)
      11'b00000000000 : romData <= 32'hEFBEADDE;
      11'b00000000001 : romData <= 32'h00000015;
      11'b00000000010 : romData <= 32'h11000000;
      11'b00000000011 : romData <= 32'h00000015;
      11'b00000000100 : romData <= 32'h0F000000;
      11'b00000000101 : romData <= 32'h00000015;
      11'b00000000110 : romData <= 32'h0D000000;
      11'b00000000111 : romData <= 32'h00000015;
      11'b00000001000 : romData <= 32'h0B000000;
      11'b00000001001 : romData <= 32'h00000015;
      11'b00000001010 : romData <= 32'h09000000;
      11'b00000001011 : romData <= 32'h00000015;
      11'b00000001100 : romData <= 32'h00C02018;
      11'b00000001101 : romData <= 32'hFC1F21A8;
      11'b00000001110 : romData <= 32'h050060E0;
      11'b00000001111 : romData <= 32'hF3020004;
      11'b00000010000 : romData <= 32'h050080E0;
      11'b00000010010 : romData <= 32'h00000015;
      11'b00000010011 : romData <= 32'h84FF219C;
      11'b00000010100 : romData <= 32'h001001D4;
      11'b00000010101 : romData <= 32'h041801D4;
      11'b00000010110 : romData <= 32'h082001D4;
      11'b00000010111 : romData <= 32'h0C2801D4;
      11'b00000011000 : romData <= 32'h103001D4;
      11'b00000011001 : romData <= 32'h143801D4;
      11'b00000011010 : romData <= 32'h184001D4;
      11'b00000011011 : romData <= 32'h1C4801D4;
      11'b00000011100 : romData <= 32'h205001D4;
      11'b00000011101 : romData <= 32'h245801D4;
      11'b00000011110 : romData <= 32'h286001D4;
      11'b00000011111 : romData <= 32'h2C6801D4;
      11'b00000100000 : romData <= 32'h307001D4;
      11'b00000100001 : romData <= 32'h347801D4;
      11'b00000100010 : romData <= 32'h388001D4;
      11'b00000100011 : romData <= 32'h3C8801D4;
      11'b00000100100 : romData <= 32'h409001D4;
      11'b00000100101 : romData <= 32'h449801D4;
      11'b00000100110 : romData <= 32'h48A001D4;
      11'b00000100111 : romData <= 32'h4CA801D4;
      11'b00000101000 : romData <= 32'h50B001D4;
      11'b00000101001 : romData <= 32'h54B801D4;
      11'b00000101010 : romData <= 32'h58C001D4;
      11'b00000101011 : romData <= 32'h5CC801D4;
      11'b00000101100 : romData <= 32'h60D001D4;
      11'b00000101101 : romData <= 32'h64D801D4;
      11'b00000101110 : romData <= 32'h68E001D4;
      11'b00000101111 : romData <= 32'h6CE801D4;
      11'b00000110000 : romData <= 32'h70F001D4;
      11'b00000110001 : romData <= 32'h74F801D4;
      11'b00000110010 : romData <= 32'h1200E0B7;
      11'b00000110011 : romData <= 32'h0200FFBB;
      11'b00000110100 : romData <= 32'h00F0C01B;
      11'b00000110101 : romData <= 32'h6C01DEAB;
      11'b00000110110 : romData <= 32'h00F8DEE3;
      11'b00000110111 : romData <= 32'h0000FE87;
      11'b00000111000 : romData <= 32'h00F80048;
      11'b00000111001 : romData <= 32'h00000015;
      11'b00000111010 : romData <= 32'h00004184;
      11'b00000111011 : romData <= 32'h04006184;
      11'b00000111100 : romData <= 32'h08008184;
      11'b00000111101 : romData <= 32'h0C00A184;
      11'b00000111110 : romData <= 32'h1000C184;
      11'b00000111111 : romData <= 32'h1400E184;
      11'b00001000000 : romData <= 32'h18000185;
      11'b00001000001 : romData <= 32'h1C002185;
      11'b00001000010 : romData <= 32'h20004185;
      11'b00001000011 : romData <= 32'h24006185;
      11'b00001000100 : romData <= 32'h28008185;
      11'b00001000101 : romData <= 32'h2C00A185;
      11'b00001000110 : romData <= 32'h3000C185;
      11'b00001000111 : romData <= 32'h3400E185;
      11'b00001001000 : romData <= 32'h38000186;
      11'b00001001001 : romData <= 32'h3C002186;
      11'b00001001010 : romData <= 32'h40004186;
      11'b00001001011 : romData <= 32'h44006186;
      11'b00001001100 : romData <= 32'h48008186;
      11'b00001001101 : romData <= 32'h4C00A186;
      11'b00001001110 : romData <= 32'h5000C186;
      11'b00001001111 : romData <= 32'h5400E186;
      11'b00001010000 : romData <= 32'h58000187;
      11'b00001010001 : romData <= 32'h5C002187;
      11'b00001010010 : romData <= 32'h60004187;
      11'b00001010011 : romData <= 32'h64006187;
      11'b00001010100 : romData <= 32'h68008187;
      11'b00001010101 : romData <= 32'h6C00A187;
      11'b00001010110 : romData <= 32'h7000C187;
      11'b00001010111 : romData <= 32'h7400E187;
      11'b00001011000 : romData <= 32'h7C00219C;
      11'b00001011001 : romData <= 32'h00000024;
      11'b00001011010 : romData <= 32'h00000015;
      11'b00001011011 : romData <= 32'h300000F0;
      11'b00001011100 : romData <= 32'h840100F0;
      11'b00001011101 : romData <= 32'hA00100F0;
      11'b00001011110 : romData <= 32'hBC0100F0;
      11'b00001011111 : romData <= 32'hD80100F0;
      11'b00001100000 : romData <= 32'hF40100F0;
      11'b00001100001 : romData <= 32'h00F0A018;
      11'b00001100010 : romData <= 32'h00F08018;
      11'b00001100011 : romData <= 32'h00F06018;
      11'b00001100100 : romData <= 32'hC017A59C;
      11'b00001100101 : romData <= 32'h8C08849C;
      11'b00001100110 : romData <= 32'h39010000;
      11'b00001100111 : romData <= 32'hF409639C;
      11'b00001101000 : romData <= 32'h00F0A018;
      11'b00001101001 : romData <= 32'h00F08018;
      11'b00001101010 : romData <= 32'h00F06018;
      11'b00001101011 : romData <= 32'hCB17A59C;
      11'b00001101100 : romData <= 32'h8C08849C;
      11'b00001101101 : romData <= 32'h32010000;
      11'b00001101110 : romData <= 32'hF409639C;
      11'b00001101111 : romData <= 32'h00F0A018;
      11'b00001110000 : romData <= 32'h00F08018;
      11'b00001110001 : romData <= 32'h00F06018;
      11'b00001110010 : romData <= 32'hD517A59C;
      11'b00001110011 : romData <= 32'h8C08849C;
      11'b00001110100 : romData <= 32'h2B010000;
      11'b00001110101 : romData <= 32'hF409639C;
      11'b00001110110 : romData <= 32'h00F0A018;
      11'b00001110111 : romData <= 32'h00F08018;
      11'b00001111000 : romData <= 32'h00F06018;
      11'b00001111001 : romData <= 32'hDA17A59C;
      11'b00001111010 : romData <= 32'h8C08849C;
      11'b00001111011 : romData <= 32'h24010000;
      11'b00001111100 : romData <= 32'hF409639C;
      11'b00001111101 : romData <= 32'h00F0A018;
      11'b00001111110 : romData <= 32'h00F08018;
      11'b00001111111 : romData <= 32'h00F06018;
      11'b00010000000 : romData <= 32'hDF17A59C;
      11'b00010000001 : romData <= 32'h8C08849C;
      11'b00010000010 : romData <= 32'h1D010000;
      11'b00010000011 : romData <= 32'hF409639C;
      11'b00010000100 : romData <= 32'h0000601A;
      11'b00010000101 : romData <= 32'h0700A0AA;
      11'b00010000110 : romData <= 32'h02A83372;
      11'b00010000111 : romData <= 32'h0000E01A;
      11'b00010001000 : romData <= 32'h010031A6;
      11'b00010001001 : romData <= 32'h00B831E4;
      11'b00010001010 : romData <= 32'hFCFFFF13;
      11'b00010001011 : romData <= 32'h00000015;
      11'b00010001100 : romData <= 32'h00480044;
      11'b00010001101 : romData <= 32'h00000015;
      11'b00010001110 : romData <= 32'h00006019;
      11'b00010001111 : romData <= 32'h02186B71;
      11'b00010010000 : romData <= 32'h00480044;
      11'b00010010001 : romData <= 32'h00000015;
      11'b00010010010 : romData <= 32'h160020AA;
      11'b00010010011 : romData <= 32'h02890370;
      11'b00010010100 : romData <= 32'h020020AA;
      11'b00010010101 : romData <= 32'h070060AA;
      11'b00010010110 : romData <= 32'h02991170;
      11'b00010010111 : romData <= 32'hEDFFFF03;
      11'b00010011000 : romData <= 32'h00000015;
      11'b00010011001 : romData <= 32'hDCFF219C;
      11'b00010011010 : romData <= 32'h008001D4;
      11'b00010011011 : romData <= 32'h049001D4;
      11'b00010011100 : romData <= 32'h08A001D4;
      11'b00010011101 : romData <= 32'h0CB001D4;
      11'b00010011110 : romData <= 32'h10C001D4;
      11'b00010011111 : romData <= 32'h14D001D4;
      11'b00010100000 : romData <= 32'h18E001D4;
      11'b00010100001 : romData <= 32'h1CF001D4;
      11'b00010100010 : romData <= 32'h204801D4;
      11'b00010100011 : romData <= 32'h0418C3E2;
      11'b00010100100 : romData <= 32'h042044E2;
      11'b00010100101 : romData <= 32'h0000001A;
      11'b00010100110 : romData <= 32'h0000801A;
      11'b00010100111 : romData <= 32'h160000AB;
      11'b00010101000 : romData <= 32'h200040AB;
      11'b00010101001 : romData <= 32'h010080AB;
      11'b00010101010 : romData <= 32'h0700C0AB;
      11'b00010101011 : romData <= 32'h009094E5;
      11'b00010101100 : romData <= 32'h0C000010;
      11'b00010101101 : romData <= 32'h20002185;
      11'b00010101110 : romData <= 32'h00000186;
      11'b00010101111 : romData <= 32'h04004186;
      11'b00010110000 : romData <= 32'h08008186;
      11'b00010110001 : romData <= 32'h0C00C186;
      11'b00010110010 : romData <= 32'h10000187;
      11'b00010110011 : romData <= 32'h14004187;
      11'b00010110100 : romData <= 32'h18008187;
      11'b00010110101 : romData <= 32'h1C00C187;
      11'b00010110110 : romData <= 32'h00480044;
      11'b00010110111 : romData <= 32'h2400219C;
      11'b00010111000 : romData <= 32'h02C11070;
      11'b00010111001 : romData <= 32'h180020AA;
      11'b00010111010 : romData <= 32'h008076E2;
      11'b00010111011 : romData <= 32'h0000B386;
      11'b00010111100 : romData <= 32'h0102B572;
      11'b00010111101 : romData <= 32'h02891570;
      11'b00010111110 : romData <= 32'h0100319E;
      11'b00010111111 : romData <= 32'h00D031E4;
      11'b00011000000 : romData <= 32'hFBFFFF13;
      11'b00011000001 : romData <= 32'h0400739E;
      11'b00011000010 : romData <= 32'h02F11C70;
      11'b00011000011 : romData <= 32'hC1FFFF07;
      11'b00011000100 : romData <= 32'h0800949E;
      11'b00011000101 : romData <= 32'hE6FFFF03;
      11'b00011000110 : romData <= 32'h2000109E;
      11'b00011000111 : romData <= 32'hB4FF219C;
      11'b00011001000 : romData <= 32'h00F08018;
      11'b00011001001 : romData <= 32'h2000A0A8;
      11'b00011001010 : romData <= 32'h7C1E849C;
      11'b00011001011 : romData <= 32'h0C00619C;
      11'b00011001100 : romData <= 32'h2C8001D4;
      11'b00011001101 : romData <= 32'h309001D4;
      11'b00011001110 : romData <= 32'h38B001D4;
      11'b00011001111 : romData <= 32'h3CC001D4;
      11'b00011010000 : romData <= 32'h40D001D4;
      11'b00011010001 : romData <= 32'h44E001D4;
      11'b00011010010 : romData <= 32'h484801D4;
      11'b00011010011 : romData <= 32'h34A001D4;
      11'b00011010100 : romData <= 32'hAE010004;
      11'b00011010101 : romData <= 32'h00F0401A;
      11'b00011010110 : romData <= 32'h00F0001A;
      11'b00011010111 : romData <= 32'h8C08529E;
      11'b00011011000 : romData <= 32'hF409109E;
      11'b00011011001 : romData <= 32'h00F0A018;
      11'b00011011010 : romData <= 32'hE817A59C;
      11'b00011011011 : romData <= 32'h049092E0;
      11'b00011011100 : romData <= 32'hC3000004;
      11'b00011011101 : romData <= 32'h048070E0;
      11'b00011011110 : romData <= 32'h1F00201A;
      11'b00011011111 : romData <= 32'h00F0C01A;
      11'b00011100000 : romData <= 32'h0000601A;
      11'b00011100001 : romData <= 32'h00FC31AA;
      11'b00011100010 : romData <= 32'h0004001B;
      11'b00011100011 : romData <= 32'hFFFF40AF;
      11'b00011100100 : romData <= 32'h1918D69E;
      11'b00011100101 : romData <= 32'h010080AB;
      11'b00011100110 : romData <= 32'h0200A0AA;
      11'b00011100111 : romData <= 32'h08A891E2;
      11'b00011101000 : romData <= 32'h00C094E2;
      11'b00011101001 : romData <= 32'h0000B486;
      11'b00011101010 : romData <= 32'h00D015E4;
      11'b00011101011 : romData <= 32'h1D000010;
      11'b00011101100 : romData <= 32'h0100319E;
      11'b00011101101 : romData <= 32'h0000201A;
      11'b00011101110 : romData <= 32'h008813E4;
      11'b00011101111 : romData <= 32'h10000010;
      11'b00011110000 : romData <= 32'h04B0B6E0;
      11'b00011110001 : romData <= 32'h00F0A018;
      11'b00011110010 : romData <= 32'h0B18A59C;
      11'b00011110011 : romData <= 32'h049092E0;
      11'b00011110100 : romData <= 32'h048070E0;
      11'b00011110101 : romData <= 32'h30004186;
      11'b00011110110 : romData <= 32'h2C000186;
      11'b00011110111 : romData <= 32'h34008186;
      11'b00011111000 : romData <= 32'h3800C186;
      11'b00011111001 : romData <= 32'h3C000187;
      11'b00011111010 : romData <= 32'h40004187;
      11'b00011111011 : romData <= 32'h44008187;
      11'b00011111100 : romData <= 32'h48002185;
      11'b00011111101 : romData <= 32'hA2000000;
      11'b00011111110 : romData <= 32'h4C00219C;
      11'b00011111111 : romData <= 32'h049092E0;
      11'b00100000000 : romData <= 32'h9F000004;
      11'b00100000001 : romData <= 32'h048070E0;
      11'b00100000010 : romData <= 32'h90FFFF07;
      11'b00100000011 : romData <= 32'h04A074E0;
      11'b00100000100 : romData <= 32'h1F00201A;
      11'b00100000101 : romData <= 32'h04E07CE2;
      11'b00100000110 : romData <= 32'h00FC31AA;
      11'b00100000111 : romData <= 32'h0100319E;
      11'b00100001000 : romData <= 32'h2000A01A;
      11'b00100001001 : romData <= 32'h00A831E4;
      11'b00100001010 : romData <= 32'hDDFFFF13;
      11'b00100001011 : romData <= 32'h0200A0AA;
      11'b00100001100 : romData <= 32'h00F0A018;
      11'b00100001101 : romData <= 32'h3518A59C;
      11'b00100001110 : romData <= 32'h049092E0;
      11'b00100001111 : romData <= 32'h90000004;
      11'b00100010000 : romData <= 32'h048070E0;
      11'b00100010001 : romData <= 32'h0C00819E;
      11'b00100010010 : romData <= 32'h04A074E2;
      11'b00100010011 : romData <= 32'h180020AA;
      11'b00100010100 : romData <= 32'h2000E0AA;
      11'b00100010101 : romData <= 32'h0000B386;
      11'b00100010110 : romData <= 32'h0102B572;
      11'b00100010111 : romData <= 32'h02891570;
      11'b00100011000 : romData <= 32'h0100319E;
      11'b00100011001 : romData <= 32'h00B831E4;
      11'b00100011010 : romData <= 32'hFBFFFF13;
      11'b00100011011 : romData <= 32'h0400739E;
      11'b00100011100 : romData <= 32'h7F00201A;
      11'b00100011101 : romData <= 32'h00F031AA;
      11'b00100011110 : romData <= 32'h160060AA;
      11'b00100011111 : romData <= 32'h02991170;
      11'b00100100000 : romData <= 32'h010020AA;
      11'b00100100001 : romData <= 32'h070060AA;
      11'b00100100010 : romData <= 32'h02991170;
      11'b00100100011 : romData <= 32'h61FFFF07;
      11'b00100100100 : romData <= 32'h00000015;
      11'b00100100101 : romData <= 32'h00F0A018;
      11'b00100100110 : romData <= 32'h5618A59C;
      11'b00100100111 : romData <= 32'h049092E0;
      11'b00100101000 : romData <= 32'h77000004;
      11'b00100101001 : romData <= 32'h048070E0;
      11'b00100101010 : romData <= 32'h7F04201A;
      11'b00100101011 : romData <= 32'h00F031AA;
      11'b00100101100 : romData <= 32'h0000601A;
      11'b00100101101 : romData <= 32'h080020AB;
      11'b00100101110 : romData <= 32'h0000B186;
      11'b00100101111 : romData <= 32'h0000F486;
      11'b00100110000 : romData <= 32'h00A817E4;
      11'b00100110001 : romData <= 32'h14000010;
      11'b00100110010 : romData <= 32'h0400319E;
      11'b00100110011 : romData <= 32'h00F0A018;
      11'b00100110100 : romData <= 32'h08B801D4;
      11'b00100110101 : romData <= 32'h04A801D4;
      11'b00100110110 : romData <= 32'h009801D4;
      11'b00100110111 : romData <= 32'h049092E0;
      11'b00100111000 : romData <= 32'h048070E0;
      11'b00100111001 : romData <= 32'h66000004;
      11'b00100111010 : romData <= 32'h7B18A59C;
      11'b00100111011 : romData <= 32'h48002185;
      11'b00100111100 : romData <= 32'h2C000186;
      11'b00100111101 : romData <= 32'h30004186;
      11'b00100111110 : romData <= 32'h34008186;
      11'b00100111111 : romData <= 32'h3800C186;
      11'b00101000000 : romData <= 32'h3C000187;
      11'b00101000001 : romData <= 32'h40004187;
      11'b00101000010 : romData <= 32'h44008187;
      11'b00101000011 : romData <= 32'h00480044;
      11'b00101000100 : romData <= 32'h4C00219C;
      11'b00101000101 : romData <= 32'h0100739E;
      11'b00101000110 : romData <= 32'h00C833E4;
      11'b00101000111 : romData <= 32'hE7FFFF13;
      11'b00101001000 : romData <= 32'h0400949E;
      11'b00101001001 : romData <= 32'h00F0A018;
      11'b00101001010 : romData <= 32'hA9FFFF03;
      11'b00101001011 : romData <= 32'h9B18A59C;
      11'b00101001100 : romData <= 32'hE8FF219C;
      11'b00101001101 : romData <= 32'h008001D4;
      11'b00101001110 : romData <= 32'h049001D4;
      11'b00101001111 : romData <= 32'h08A001D4;
      11'b00101010000 : romData <= 32'h0CB001D4;
      11'b00101010001 : romData <= 32'h10C001D4;
      11'b00101010010 : romData <= 32'h144801D4;
      11'b00101010011 : romData <= 32'h041843E2;
      11'b00101010100 : romData <= 32'h042084E2;
      11'b00101010101 : romData <= 32'h1C0000AA;
      11'b00101010110 : romData <= 32'h090000AB;
      11'b00101010111 : romData <= 32'hFCFFC0AE;
      11'b00101011000 : romData <= 32'h488074E0;
      11'b00101011001 : romData <= 32'h0F0023A6;
      11'b00101011010 : romData <= 32'h00C051E4;
      11'b00101011011 : romData <= 32'h03000010;
      11'b00101011100 : romData <= 32'h3700719C;
      11'b00101011101 : romData <= 32'h3000719C;
      11'b00101011110 : romData <= 32'h00900048;
      11'b00101011111 : romData <= 32'hFCFF109E;
      11'b00101100000 : romData <= 32'h00B030E4;
      11'b00101100001 : romData <= 32'hF8FFFF13;
      11'b00101100010 : romData <= 32'h488074E0;
      11'b00101100011 : romData <= 32'h00000186;
      11'b00101100100 : romData <= 32'h04004186;
      11'b00101100101 : romData <= 32'h08008186;
      11'b00101100110 : romData <= 32'h0C00C186;
      11'b00101100111 : romData <= 32'h10000187;
      11'b00101101000 : romData <= 32'h14002185;
      11'b00101101001 : romData <= 32'h00480044;
      11'b00101101010 : romData <= 32'h1800219C;
      11'b00101101011 : romData <= 32'hDCFF219C;
      11'b00101101100 : romData <= 32'h0C8001D4;
      11'b00101101101 : romData <= 32'h109001D4;
      11'b00101101110 : romData <= 32'h14A001D4;
      11'b00101101111 : romData <= 32'h18B001D4;
      11'b00101110000 : romData <= 32'h1CC001D4;
      11'b00101110001 : romData <= 32'h204801D4;
      11'b00101110010 : romData <= 32'h0418C3E2;
      11'b00101110011 : romData <= 32'h042044E2;
      11'b00101110100 : romData <= 32'h0000801A;
      11'b00101110101 : romData <= 32'h0000001A;
      11'b00101110110 : romData <= 32'h0A0000AB;
      11'b00101110111 : romData <= 32'h04C098E0;
      11'b00101111000 : romData <= 32'h73040004;
      11'b00101111001 : romData <= 32'h049072E0;
      11'b00101111010 : romData <= 32'h0200219E;
      11'b00101111011 : romData <= 32'h00A031E2;
      11'b00101111100 : romData <= 32'h30006B9D;
      11'b00101111101 : romData <= 32'h005811D8;
      11'b00101111110 : romData <= 32'h0000201A;
      11'b00101111111 : romData <= 32'h008814E4;
      11'b00110000000 : romData <= 32'h04000010;
      11'b00110000001 : romData <= 32'h008812E4;
      11'b00110000010 : romData <= 32'h05000010;
      11'b00110000011 : romData <= 32'h049072E0;
      11'b00110000100 : romData <= 32'h0100109E;
      11'b00110000101 : romData <= 32'hFF0010A6;
      11'b00110000110 : romData <= 32'h049072E0;
      11'b00110000111 : romData <= 32'h4B040004;
      11'b00110001000 : romData <= 32'h04C098E0;
      11'b00110001001 : romData <= 32'h0100949E;
      11'b00110001010 : romData <= 32'h00C034E4;
      11'b00110001011 : romData <= 32'hECFFFF13;
      11'b00110001100 : romData <= 32'h04584BE2;
      11'b00110001101 : romData <= 32'h0000201A;
      11'b00110001110 : romData <= 32'h008830E4;
      11'b00110001111 : romData <= 32'h0A000010;
      11'b00110010000 : romData <= 32'hFFFF109E;
      11'b00110010001 : romData <= 32'h0C000186;
      11'b00110010010 : romData <= 32'h10004186;
      11'b00110010011 : romData <= 32'h14008186;
      11'b00110010100 : romData <= 32'h1800C186;
      11'b00110010101 : romData <= 32'h1C000187;
      11'b00110010110 : romData <= 32'h20002185;
      11'b00110010111 : romData <= 32'h00480044;
      11'b00110011000 : romData <= 32'h2400219C;
      11'b00110011001 : romData <= 32'h0200219E;
      11'b00110011010 : romData <= 32'h008031E2;
      11'b00110011011 : romData <= 32'h00B00048;
      11'b00110011100 : romData <= 32'h0000718C;
      11'b00110011101 : romData <= 32'hF1FFFF03;
      11'b00110011110 : romData <= 32'h0000201A;
      11'b00110011111 : romData <= 32'hE0FF219C;
      11'b00110100000 : romData <= 32'h008001D4;
      11'b00110100001 : romData <= 32'h049001D4;
      11'b00110100010 : romData <= 32'h08A001D4;
      11'b00110100011 : romData <= 32'h0CB001D4;
      11'b00110100100 : romData <= 32'h14D001D4;
      11'b00110100101 : romData <= 32'h18E001D4;
      11'b00110100110 : romData <= 32'h10C001D4;
      11'b00110100111 : romData <= 32'h1C4801D4;
      11'b00110101000 : romData <= 32'h041883E2;
      11'b00110101001 : romData <= 32'h042004E2;
      11'b00110101010 : romData <= 32'h042845E2;
      11'b00110101011 : romData <= 32'h2000C19E;
      11'b00110101100 : romData <= 32'h250040AB;
      11'b00110101101 : romData <= 32'h630080AB;
      11'b00110101110 : romData <= 32'h00007290;
      11'b00110101111 : romData <= 32'h0000201A;
      11'b00110110000 : romData <= 32'h008823E4;
      11'b00110110001 : romData <= 32'h3B00000C;
      11'b00110110010 : romData <= 32'h00D023E4;
      11'b00110110011 : romData <= 32'h5A000010;
      11'b00110110100 : romData <= 32'hFF0003A7;
      11'b00110110101 : romData <= 32'h01003292;
      11'b00110110110 : romData <= 32'h00E011E4;
      11'b00110110111 : romData <= 32'h4D000010;
      11'b00110111000 : romData <= 32'h00E051E5;
      11'b00110111001 : romData <= 32'h1B000010;
      11'b00110111010 : romData <= 32'h0000601A;
      11'b00110111011 : romData <= 32'h009811E4;
      11'b00110111100 : romData <= 32'h28000010;
      11'b00110111101 : romData <= 32'h580060AA;
      11'b00110111110 : romData <= 32'h009811E4;
      11'b00110111111 : romData <= 32'h37000010;
      11'b00111000000 : romData <= 32'h0400169F;
      11'b00111000001 : romData <= 32'h00A00048;
      11'b00111000010 : romData <= 32'h250060A8;
      11'b00111000011 : romData <= 32'h0000201A;
      11'b00111000100 : romData <= 32'h008810E4;
      11'b00111000101 : romData <= 32'h04000010;
      11'b00111000110 : romData <= 32'h00000015;
      11'b00111000111 : romData <= 32'h00800048;
      11'b00111001000 : romData <= 32'h250060A8;
      11'b00111001001 : romData <= 32'h0100128F;
      11'b00111001010 : romData <= 32'h00A00048;
      11'b00111001011 : romData <= 32'h04C078E0;
      11'b00111001100 : romData <= 32'h0000201A;
      11'b00111001101 : romData <= 32'h008810E4;
      11'b00111001110 : romData <= 32'h33000010;
      11'b00111001111 : romData <= 32'h00000015;
      11'b00111010000 : romData <= 32'h00800048;
      11'b00111010001 : romData <= 32'h04C078E0;
      11'b00111010010 : romData <= 32'h30000000;
      11'b00111010011 : romData <= 32'h0100529E;
      11'b00111010100 : romData <= 32'h640060AA;
      11'b00111010101 : romData <= 32'h009811E4;
      11'b00111010110 : romData <= 32'hEBFFFF0F;
      11'b00111010111 : romData <= 32'h0400169F;
      11'b00111011000 : romData <= 32'h04A074E0;
      11'b00111011001 : romData <= 32'h0000D686;
      11'b00111011010 : romData <= 32'h91FFFF07;
      11'b00111011011 : romData <= 32'h04B096E0;
      11'b00111011100 : romData <= 32'h0000201A;
      11'b00111011101 : romData <= 32'h008810E4;
      11'b00111011110 : romData <= 32'h22000010;
      11'b00111011111 : romData <= 32'h04B096E0;
      11'b00111100000 : romData <= 32'h8BFFFF07;
      11'b00111100001 : romData <= 32'h048070E0;
      11'b00111100010 : romData <= 32'h1F000000;
      11'b00111100011 : romData <= 32'h04C0D8E2;
      11'b00111100100 : romData <= 32'h00A00048;
      11'b00111100101 : romData <= 32'h04D07AE0;
      11'b00111100110 : romData <= 32'h0000201A;
      11'b00111100111 : romData <= 32'h008810E4;
      11'b00111101000 : romData <= 32'h04000010;
      11'b00111101001 : romData <= 32'h04D07AE0;
      11'b00111101010 : romData <= 32'h00800048;
      11'b00111101011 : romData <= 32'h00000015;
      11'b00111101100 : romData <= 32'h00000186;
      11'b00111101101 : romData <= 32'h04004186;
      11'b00111101110 : romData <= 32'h08008186;
      11'b00111101111 : romData <= 32'h0C00C186;
      11'b00111110000 : romData <= 32'h10000187;
      11'b00111110001 : romData <= 32'h14004187;
      11'b00111110010 : romData <= 32'h18008187;
      11'b00111110011 : romData <= 32'h1C002185;
      11'b00111110100 : romData <= 32'h00480044;
      11'b00111110101 : romData <= 32'h2000219C;
      11'b00111110110 : romData <= 32'h04A074E0;
      11'b00111110111 : romData <= 32'h0000D686;
      11'b00111111000 : romData <= 32'h54FFFF07;
      11'b00111111001 : romData <= 32'h04B096E0;
      11'b00111111010 : romData <= 32'h0000201A;
      11'b00111111011 : romData <= 32'h008810E4;
      11'b00111111100 : romData <= 32'h04000010;
      11'b00111111101 : romData <= 32'h04B096E0;
      11'b00111111110 : romData <= 32'h4EFFFF07;
      11'b00111111111 : romData <= 32'h048070E0;
      11'b01000000000 : romData <= 32'h04C0D8E2;
      11'b01000000001 : romData <= 32'h0100529E;
      11'b01000000010 : romData <= 32'hACFFFF03;
      11'b01000000011 : romData <= 32'h0100529E;
      11'b01000000100 : romData <= 32'h0300568E;
      11'b01000000101 : romData <= 32'h00A00048;
      11'b01000000110 : romData <= 32'h049072E0;
      11'b01000000111 : romData <= 32'h0000201A;
      11'b01000001000 : romData <= 32'h008810E4;
      11'b01000001001 : romData <= 32'hE3FFFF13;
      11'b01000001010 : romData <= 32'h049072E0;
      11'b01000001011 : romData <= 32'hDFFFFF03;
      11'b01000001100 : romData <= 32'h00000015;
      11'b01000001101 : romData <= 32'h00A00048;
      11'b01000001110 : romData <= 32'h04C078E0;
      11'b01000001111 : romData <= 32'h0000201A;
      11'b01000010000 : romData <= 32'h008810E4;
      11'b01000010001 : romData <= 32'hF1FFFF13;
      11'b01000010010 : romData <= 32'h00000015;
      11'b01000010011 : romData <= 32'h00800048;
      11'b01000010100 : romData <= 32'h04C078E0;
      11'b01000010101 : romData <= 32'h99FFFF03;
      11'b01000010110 : romData <= 32'h0100529E;
      11'b01000010111 : romData <= 32'h0050201A;
      11'b01000011000 : romData <= 32'h030071AA;
      11'b01000011001 : romData <= 32'h83FFA0AE;
      11'b01000011010 : romData <= 32'h00A813D8;
      11'b01000011011 : romData <= 32'h2800A0AA;
      11'b01000011100 : romData <= 32'h00A811D8;
      11'b01000011101 : romData <= 32'h010031AA;
      11'b01000011110 : romData <= 32'h000011D8;
      11'b01000011111 : romData <= 32'h030020AA;
      11'b01000100000 : romData <= 32'h008813D8;
      11'b01000100001 : romData <= 32'h00480044;
      11'b01000100010 : romData <= 32'h00000015;
      11'b01000100011 : romData <= 32'h0050601A;
      11'b01000100100 : romData <= 32'hFF0063A4;
      11'b01000100101 : romData <= 32'h0500B3AA;
      11'b01000100110 : romData <= 32'h0000358E;
      11'b01000100111 : romData <= 32'h400031A6;
      11'b01000101000 : romData <= 32'h0000E01A;
      11'b01000101001 : romData <= 32'h00B811E4;
      11'b01000101010 : romData <= 32'h05000010;
      11'b01000101011 : romData <= 32'h00000015;
      11'b01000101100 : romData <= 32'h001813D8;
      11'b01000101101 : romData <= 32'h00480044;
      11'b01000101110 : romData <= 32'h00000015;
      11'b01000101111 : romData <= 32'h00000015;
      11'b01000110000 : romData <= 32'hF6FFFF03;
      11'b01000110001 : romData <= 32'h00000015;
      11'b01000110010 : romData <= 32'h0050601A;
      11'b01000110011 : romData <= 32'h0500B3AA;
      11'b01000110100 : romData <= 32'h0000358E;
      11'b01000110101 : romData <= 32'h010031A6;
      11'b01000110110 : romData <= 32'h0000E01A;
      11'b01000110111 : romData <= 32'h00B811E4;
      11'b01000111000 : romData <= 32'hFCFFFF13;
      11'b01000111001 : romData <= 32'h00000015;
      11'b01000111010 : romData <= 32'h0000738D;
      11'b01000111011 : romData <= 32'h00480044;
      11'b01000111100 : romData <= 32'h00000015;
      11'b01000111101 : romData <= 32'hF0FF219C;
      11'b01000111110 : romData <= 32'hFF0063A4;
      11'b01000111111 : romData <= 32'h008001D4;
      11'b01001000000 : romData <= 32'hD0FF039E;
      11'b01001000001 : romData <= 32'hFF0030A6;
      11'b01001000010 : romData <= 32'h090060AA;
      11'b01001000011 : romData <= 32'h049001D4;
      11'b01001000100 : romData <= 32'h08A001D4;
      11'b01001000101 : romData <= 32'h009851E4;
      11'b01001000110 : romData <= 32'h0800000C;
      11'b01001000111 : romData <= 32'h0C4801D4;
      11'b01001001000 : romData <= 32'hBFFF239E;
      11'b01001001001 : romData <= 32'hFF0031A6;
      11'b01001001010 : romData <= 32'h050060AA;
      11'b01001001011 : romData <= 32'h009851E4;
      11'b01001001100 : romData <= 32'h18000010;
      11'b01001001101 : romData <= 32'hC9FF039E;
      11'b01001001110 : romData <= 32'h090040AA;
      11'b01001001111 : romData <= 32'h050080AA;
      11'b01001010000 : romData <= 32'hE2FFFF07;
      11'b01001010001 : romData <= 32'h00000015;
      11'b01001010010 : romData <= 32'hFF006BA5;
      11'b01001010011 : romData <= 32'hD0FF2B9E;
      11'b01001010100 : romData <= 32'hFF0071A6;
      11'b01001010101 : romData <= 32'h009053E4;
      11'b01001010110 : romData <= 32'h04000010;
      11'b01001010111 : romData <= 32'h0400A0AA;
      11'b01001011000 : romData <= 32'h08A810E2;
      11'b01001011001 : romData <= 32'h008011E2;
      11'b01001011010 : romData <= 32'hBFFF2B9E;
      11'b01001011011 : romData <= 32'hFF0031A6;
      11'b01001011100 : romData <= 32'h00A051E4;
      11'b01001011101 : romData <= 32'h10000010;
      11'b01001011110 : romData <= 32'h9FFF2B9E;
      11'b01001011111 : romData <= 32'h040020AA;
      11'b01001100000 : romData <= 32'h088810E2;
      11'b01001100001 : romData <= 32'hC9FF6B9D;
      11'b01001100010 : romData <= 32'hEEFFFF03;
      11'b01001100011 : romData <= 32'h00800BE2;
      11'b01001100100 : romData <= 32'h9FFF239E;
      11'b01001100101 : romData <= 32'hFF0031A6;
      11'b01001100110 : romData <= 32'h009851E4;
      11'b01001100111 : romData <= 32'h04000010;
      11'b01001101000 : romData <= 32'h00000015;
      11'b01001101001 : romData <= 32'hE5FFFF03;
      11'b01001101010 : romData <= 32'hA9FF039E;
      11'b01001101011 : romData <= 32'hE3FFFF03;
      11'b01001101100 : romData <= 32'h0000001A;
      11'b01001101101 : romData <= 32'hFF0031A6;
      11'b01001101110 : romData <= 32'h00A051E4;
      11'b01001101111 : romData <= 32'h05000010;
      11'b01001110000 : romData <= 32'h040020AA;
      11'b01001110001 : romData <= 32'h088810E2;
      11'b01001110010 : romData <= 32'hF0FFFF03;
      11'b01001110011 : romData <= 32'hA9FF6B9D;
      11'b01001110100 : romData <= 32'h0090B3E4;
      11'b01001110101 : romData <= 32'hDBFFFF13;
      11'b01001110110 : romData <= 32'h048070E1;
      11'b01001110111 : romData <= 32'h04004186;
      11'b01001111000 : romData <= 32'h00000186;
      11'b01001111001 : romData <= 32'h08008186;
      11'b01001111010 : romData <= 32'h0C002185;
      11'b01001111011 : romData <= 32'h00480044;
      11'b01001111100 : romData <= 32'h1000219C;
      11'b01001111101 : romData <= 32'hFF0063A4;
      11'b01001111110 : romData <= 32'h020020AA;
      11'b01001111111 : romData <= 32'h00191170;
      11'b01010000000 : romData <= 32'h00480044;
      11'b01010000001 : romData <= 32'h00000015;
      11'b01010000010 : romData <= 32'h041863E1;
      11'b01010000011 : romData <= 32'h0000201A;
      11'b01010000100 : romData <= 32'h002831E4;
      11'b01010000101 : romData <= 32'h04000010;
      11'b01010000110 : romData <= 32'h008864E2;
      11'b01010000111 : romData <= 32'h00480044;
      11'b01010001000 : romData <= 32'h00000015;
      11'b01010001001 : romData <= 32'h0000B392;
      11'b01010001010 : romData <= 32'h00886BE2;
      11'b01010001011 : romData <= 32'h00A813D8;
      11'b01010001100 : romData <= 32'hF8FFFF03;
      11'b01010001101 : romData <= 32'h0100319E;
      11'b01010001110 : romData <= 32'hA8FF219C;
      11'b01010001111 : romData <= 32'h00F08018;
      11'b01010010000 : romData <= 32'h3800A0A8;
      11'b01010010001 : romData <= 32'h9C1E849C;
      11'b01010010010 : romData <= 32'h488001D4;
      11'b01010010011 : romData <= 32'h4C9001D4;
      11'b01010010100 : romData <= 32'h50A001D4;
      11'b01010010101 : romData <= 32'h544801D4;
      11'b01010010110 : romData <= 32'hECFFFF07;
      11'b01010010111 : romData <= 32'h1000619C;
      11'b01010011000 : romData <= 32'h030020AA;
      11'b01010011001 : romData <= 32'h00011170;
      11'b01010011010 : romData <= 32'h00F0401A;
      11'b01010011011 : romData <= 32'h00F0801A;
      11'b01010011100 : romData <= 32'h8C08529E;
      11'b01010011101 : romData <= 32'hF409949E;
      11'b01010011110 : romData <= 32'h00F0A018;
      11'b01010011111 : romData <= 32'hAE18A59C;
      11'b01010100000 : romData <= 32'h049092E0;
      11'b01010100001 : romData <= 32'hFEFEFF07;
      11'b01010100010 : romData <= 32'h04A074E0;
      11'b01010100011 : romData <= 32'h00F0A018;
      11'b01010100100 : romData <= 32'hCD18A59C;
      11'b01010100101 : romData <= 32'h049092E0;
      11'b01010100110 : romData <= 32'hF9FEFF07;
      11'b01010100111 : romData <= 32'h04A074E0;
      11'b01010101000 : romData <= 32'h00F0A018;
      11'b01010101001 : romData <= 32'hF018A59C;
      11'b01010101010 : romData <= 32'h049092E0;
      11'b01010101011 : romData <= 32'hF4FEFF07;
      11'b01010101100 : romData <= 32'h04A074E0;
      11'b01010101101 : romData <= 32'hFF00201A;
      11'b01010101110 : romData <= 32'hFFFF31AA;
      11'b01010101111 : romData <= 32'h04000072;
      11'b01010110000 : romData <= 32'h0000A01A;
      11'b01010110001 : romData <= 32'h038870E2;
      11'b01010110010 : romData <= 32'h00A813E4;
      11'b01010110011 : romData <= 32'hFCFFFF13;
      11'b01010110100 : romData <= 32'h00F0A018;
      11'b01010110101 : romData <= 32'h040020AA;
      11'b01010110110 : romData <= 32'h488830E2;
      11'b01010110111 : romData <= 32'h070031A6;
      11'b01010111000 : romData <= 32'h048801D4;
      11'b01010111001 : romData <= 32'h070030A6;
      11'b01010111010 : romData <= 32'h008801D4;
      11'b01010111011 : romData <= 32'h1D19A59C;
      11'b01010111100 : romData <= 32'h049092E0;
      11'b01010111101 : romData <= 32'hE2FEFF07;
      11'b01010111110 : romData <= 32'h04A074E0;
      11'b01010111111 : romData <= 32'h0C0020AA;
      11'b01011000000 : romData <= 32'h488830E2;
      11'b01011000001 : romData <= 32'h0F0031A6;
      11'b01011000010 : romData <= 32'h0C8801D4;
      11'b01011000011 : romData <= 32'h100020AA;
      11'b01011000100 : romData <= 32'h488830E2;
      11'b01011000101 : romData <= 32'h0F0031A6;
      11'b01011000110 : romData <= 32'h088801D4;
      11'b01011000111 : romData <= 32'h140020AA;
      11'b01011001000 : romData <= 32'h488830E2;
      11'b01011001001 : romData <= 32'h0F0031A6;
      11'b01011001010 : romData <= 32'h048801D4;
      11'b01011001011 : romData <= 32'h180020AA;
      11'b01011001100 : romData <= 32'h488830E2;
      11'b01011001101 : romData <= 32'h0F0031A6;
      11'b01011001110 : romData <= 32'h00F0A018;
      11'b01011001111 : romData <= 32'h008801D4;
      11'b01011010000 : romData <= 32'h3B19A59C;
      11'b01011010001 : romData <= 32'h049092E0;
      11'b01011010010 : romData <= 32'hCDFEFF07;
      11'b01011010011 : romData <= 32'h04A074E0;
      11'b01011010100 : romData <= 32'hADDE201A;
      11'b01011010101 : romData <= 32'h0004601A;
      11'b01011010110 : romData <= 32'hEFBE31AA;
      11'b01011010111 : romData <= 32'h0000B386;
      11'b01011011000 : romData <= 32'h008835E4;
      11'b01011011001 : romData <= 32'h13000010;
      11'b01011011010 : romData <= 32'h0000201A;
      11'b01011011011 : romData <= 32'h080010A6;
      11'b01011011100 : romData <= 32'h008830E4;
      11'b01011011101 : romData <= 32'h0F000010;
      11'b01011011110 : romData <= 32'h040033AA;
      11'b01011011111 : romData <= 32'h0200A0AA;
      11'b01011100000 : romData <= 32'h00003186;
      11'b01011100001 : romData <= 32'h08A831E2;
      11'b01011100010 : romData <= 32'h008830E4;
      11'b01011100011 : romData <= 32'h15000010;
      11'b01011100100 : romData <= 32'h0080B3E2;
      11'b01011100101 : romData <= 32'h00F0A018;
      11'b01011100110 : romData <= 32'h4C19A59C;
      11'b01011100111 : romData <= 32'h049092E0;
      11'b01011101000 : romData <= 32'hB7FEFF07;
      11'b01011101001 : romData <= 32'h04A074E0;
      11'b01011101010 : romData <= 32'h30000074;
      11'b01011101011 : romData <= 32'h00000015;
      11'b01011101100 : romData <= 32'h1000019E;
      11'b01011101101 : romData <= 32'h0000201A;
      11'b01011101110 : romData <= 32'h0000B084;
      11'b01011101111 : romData <= 32'h008825E4;
      11'b01011110000 : romData <= 32'h0D000010;
      11'b01011110001 : romData <= 32'h0400109E;
      11'b01011110010 : romData <= 32'h48000186;
      11'b01011110011 : romData <= 32'h4C004186;
      11'b01011110100 : romData <= 32'h50008186;
      11'b01011110101 : romData <= 32'h54002185;
      11'b01011110110 : romData <= 32'h00480044;
      11'b01011110111 : romData <= 32'h5800219C;
      11'b01011111000 : romData <= 32'h0000B586;
      11'b01011111001 : romData <= 32'h0400109E;
      11'b01011111010 : romData <= 32'hFCAFF0D7;
      11'b01011111011 : romData <= 32'hE8FFFF03;
      11'b01011111100 : romData <= 32'h008830E4;
      11'b01011111101 : romData <= 32'h049092E0;
      11'b01011111110 : romData <= 32'hA1FEFF07;
      11'b01011111111 : romData <= 32'h04A074E0;
      11'b01100000000 : romData <= 32'hEEFFFF03;
      11'b01100000001 : romData <= 32'h0000201A;
      11'b01100000010 : romData <= 32'hACFC219C;
      11'b01100000011 : romData <= 32'h287301D4;
      11'b01100000100 : romData <= 32'h2C8301D4;
      11'b01100000101 : romData <= 32'h309301D4;
      11'b01100000110 : romData <= 32'h44E301D4;
      11'b01100000111 : romData <= 32'h48F301D4;
      11'b01100001000 : romData <= 32'h504B01D4;
      11'b01100001001 : romData <= 32'h34A301D4;
      11'b01100001010 : romData <= 32'h38B301D4;
      11'b01100001011 : romData <= 32'h3CC301D4;
      11'b01100001100 : romData <= 32'h40D301D4;
      11'b01100001101 : romData <= 32'h0AFFFF07;
      11'b01100001110 : romData <= 32'h4C1301D4;
      11'b01100001111 : romData <= 32'h7FFFFF07;
      11'b01100010000 : romData <= 32'h010040AA;
      11'b01100010001 : romData <= 32'h00F0201A;
      11'b01100010010 : romData <= 32'h051C319E;
      11'b01100010011 : romData <= 32'h0000801B;
      11'b01100010100 : romData <= 32'h0000C019;
      11'b01100010101 : romData <= 32'h0490D2E3;
      11'b01100010110 : romData <= 32'h0000001A;
      11'b01100010111 : romData <= 32'h108801D4;
      11'b01100011000 : romData <= 32'h270040AB;
      11'b01100011001 : romData <= 32'h19FFFF07;
      11'b01100011010 : romData <= 32'h00000015;
      11'b01100011011 : romData <= 32'hFF000BA7;
      11'b01100011100 : romData <= 32'h00D018E4;
      11'b01100011101 : romData <= 32'h60020010;
      11'b01100011110 : romData <= 32'h00D058E4;
      11'b01100011111 : romData <= 32'h49000010;
      11'b01100100000 : romData <= 32'h240020AA;
      11'b01100100001 : romData <= 32'h008818E4;
      11'b01100100010 : romData <= 32'hA0000010;
      11'b01100100011 : romData <= 32'h008858E4;
      11'b01100100100 : romData <= 32'h13000010;
      11'b01100100101 : romData <= 32'h230020AA;
      11'b01100100110 : romData <= 32'h008818E4;
      11'b01100100111 : romData <= 32'h94000010;
      11'b01100101000 : romData <= 32'hF6FF789E;
      11'b01100101001 : romData <= 32'hFF0073A6;
      11'b01100101010 : romData <= 32'h160020AA;
      11'b01100101011 : romData <= 32'h008853E4;
      11'b01100101100 : romData <= 32'h09000010;
      11'b01100101101 : romData <= 32'hBFFF201A;
      11'b01100101110 : romData <= 32'hF6FF31AA;
      11'b01100101111 : romData <= 32'h889831E2;
      11'b01100110000 : romData <= 32'h010031A6;
      11'b01100110001 : romData <= 32'h0000601A;
      11'b01100110010 : romData <= 32'h009831E4;
      11'b01100110011 : romData <= 32'hE6FFFF0F;
      11'b01100110100 : romData <= 32'h00000015;
      11'b01100110101 : romData <= 32'h45000000;
      11'b01100110110 : romData <= 32'h00006019;
      11'b01100110111 : romData <= 32'h260020AA;
      11'b01100111000 : romData <= 32'h008818E4;
      11'b01100111001 : romData <= 32'hFCFFFF0F;
      11'b01100111010 : romData <= 32'h250000AB;
      11'b01100111011 : romData <= 32'hF7FEFF07;
      11'b01100111100 : romData <= 32'h0000401B;
      11'b01100111101 : romData <= 32'h00F0A018;
      11'b01100111110 : romData <= 32'h00F08018;
      11'b01100111111 : romData <= 32'h00F06018;
      11'b01101000000 : romData <= 32'h7819A59C;
      11'b01101000001 : romData <= 32'h8C08849C;
      11'b01101000010 : romData <= 32'hF409639C;
      11'b01101000011 : romData <= 32'h5CFEFF07;
      11'b01101000100 : romData <= 32'hFF004BA4;
      11'b01101000101 : romData <= 32'h200000AB;
      11'b01101000110 : romData <= 32'h00C002E4;
      11'b01101000111 : romData <= 32'h1D000010;
      11'b01101001000 : romData <= 32'h00D03AE2;
      11'b01101001001 : romData <= 32'h00D031E2;
      11'b01101001010 : romData <= 32'h2800619E;
      11'b01101001011 : romData <= 32'h0088F3E2;
      11'b01101001100 : romData <= 32'h0000A01A;
      11'b01101001101 : romData <= 32'h0100B59E;
      11'b01101001110 : romData <= 32'h001017D8;
      11'b01101001111 : romData <= 32'h188801D4;
      11'b01101010000 : romData <= 32'h14A801D4;
      11'b01101010001 : romData <= 32'hE1FEFF07;
      11'b01101010010 : romData <= 32'h0CB801D4;
      11'b01101010011 : romData <= 32'hFF004BA4;
      11'b01101010100 : romData <= 32'h00C022E4;
      11'b01101010101 : romData <= 32'h0C00E186;
      11'b01101010110 : romData <= 32'h1400A186;
      11'b01101010111 : romData <= 32'h0100F79E;
      11'b01101011000 : romData <= 32'hF5FFFF13;
      11'b01101011001 : romData <= 32'h18002186;
      11'b01101011010 : romData <= 32'h0C03319E;
      11'b01101011011 : romData <= 32'h1C00619E;
      11'b01101011100 : romData <= 32'h009831E2;
      11'b01101011101 : romData <= 32'h00A831E2;
      11'b01101011110 : romData <= 32'h0005F1DB;
      11'b01101011111 : romData <= 32'h01005A9F;
      11'b01101100000 : romData <= 32'hFF0020AA;
      11'b01101100001 : romData <= 32'h0088BAE5;
      11'b01101100010 : romData <= 32'hB6FFFF0F;
      11'b01101100011 : romData <= 32'h00000015;
      11'b01101100100 : romData <= 32'hCEFEFF07;
      11'b01101100101 : romData <= 32'h00000015;
      11'b01101100110 : romData <= 32'hE0FFFF03;
      11'b01101100111 : romData <= 32'hFF004BA4;
      11'b01101101000 : romData <= 32'h2D0020AA;
      11'b01101101001 : romData <= 32'h008818E4;
      11'b01101101010 : romData <= 32'h0B000010;
      11'b01101101011 : romData <= 32'h008858E4;
      11'b01101101100 : romData <= 32'h35000010;
      11'b01101101101 : romData <= 32'h3D0020AA;
      11'b01101101110 : romData <= 32'h2A0020AA;
      11'b01101101111 : romData <= 32'h008818E4;
      11'b01101110000 : romData <= 32'h68000010;
      11'b01101110001 : romData <= 32'h2B0020AA;
      11'b01101110010 : romData <= 32'h008818E4;
      11'b01101110011 : romData <= 32'h0700000C;
      11'b01101110100 : romData <= 32'h00006019;
      11'b01101110101 : romData <= 32'hBDFEFF07;
      11'b01101110110 : romData <= 32'h00000015;
      11'b01101110111 : romData <= 32'h180020AA;
      11'b01101111000 : romData <= 32'h08886BE1;
      11'b01101111001 : romData <= 32'h88886BE1;
      11'b01101111010 : romData <= 32'h180020AA;
      11'b01101111011 : romData <= 32'h088818E3;
      11'b01101111100 : romData <= 32'h888818E3;
      11'b01101111101 : romData <= 32'hFFFF40AC;
      11'b01101111110 : romData <= 32'h0000201A;
      11'b01101111111 : romData <= 32'hFF00E0AA;
      11'b01110000000 : romData <= 32'h008871E2;
      11'b01110000001 : romData <= 32'h008873E2;
      11'b01110000010 : romData <= 32'h0C03739E;
      11'b01110000011 : romData <= 32'h1C00A19E;
      11'b01110000100 : romData <= 32'h00A873E2;
      11'b01110000101 : romData <= 32'h00FD3393;
      11'b01110000110 : romData <= 32'h00C039E4;
      11'b01110000111 : romData <= 32'h08000010;
      11'b01110001000 : romData <= 32'h00000015;
      11'b01110001001 : romData <= 32'h01FD7392;
      11'b01110001010 : romData <= 32'h005813E4;
      11'b01110001011 : romData <= 32'h0400000C;
      11'b01110001100 : romData <= 32'h00000015;
      11'b01110001101 : romData <= 32'h048851E0;
      11'b01110001110 : romData <= 32'h000120AA;
      11'b01110001111 : romData <= 32'h0100319E;
      11'b01110010000 : romData <= 32'h00B8B1E5;
      11'b01110010001 : romData <= 32'hF0FFFF13;
      11'b01110010010 : romData <= 32'h008871E2;
      11'b01110010011 : romData <= 32'h0000201A;
      11'b01110010100 : romData <= 32'h008862E5;
      11'b01110010101 : romData <= 32'hF501000C;
      11'b01110010110 : romData <= 32'h00F0A018;
      11'b01110010111 : romData <= 32'h00F0401B;
      11'b01110011000 : romData <= 32'h00F0001B;
      11'b01110011001 : romData <= 32'h971C5A9F;
      11'b01110011010 : romData <= 32'hF409189F;
      11'b01110011011 : romData <= 32'h0000201A;
      11'b01110011100 : romData <= 32'h008832E4;
      11'b01110011101 : romData <= 32'hF0010010;
      11'b01110011110 : romData <= 32'h00881CE4;
      11'b01110011111 : romData <= 32'h79FFFF03;
      11'b01110100000 : romData <= 32'h010040AA;
      11'b01110100001 : romData <= 32'h008818E4;
      11'b01110100010 : romData <= 32'hD3FFFF13;
      11'b01110100011 : romData <= 32'h400020AA;
      11'b01110100100 : romData <= 32'h008818E4;
      11'b01110100101 : romData <= 32'hD5FFFF0F;
      11'b01110100110 : romData <= 32'h00006019;
      11'b01110100111 : romData <= 32'h96FEFF07;
      11'b01110101000 : romData <= 32'h200060A8;
      11'b01110101001 : romData <= 32'h080020AA;
      11'b01110101010 : romData <= 32'h00F0A018;
      11'b01110101011 : romData <= 32'h00F06018;
      11'b01110101100 : romData <= 32'h08888BE2;
      11'b01110101101 : romData <= 32'h005801D4;
      11'b01110101110 : romData <= 32'h0A0020AA;
      11'b01110101111 : romData <= 32'h8C19A59C;
      11'b01110110000 : romData <= 32'h00008018;
      11'b01110110001 : romData <= 32'hF409639C;
      11'b01110110010 : romData <= 32'h488894E2;
      11'b01110110011 : romData <= 32'hECFDFF07;
      11'b01110110100 : romData <= 32'h0458CBE2;
      11'b01110110101 : romData <= 32'h0000201A;
      11'b01110110110 : romData <= 32'h008814E4;
      11'b01110110111 : romData <= 32'h62FFFF0F;
      11'b01110111000 : romData <= 32'h270040AB;
      11'b01110111001 : romData <= 32'h60FFFF03;
      11'b01110111010 : romData <= 32'h0000C019;
      11'b01110111011 : romData <= 32'h00F0A018;
      11'b01110111100 : romData <= 32'h6819A59C;
      11'b01110111101 : romData <= 32'h00F08018;
      11'b01110111110 : romData <= 32'h8C08849C;
      11'b01110111111 : romData <= 32'h00F06018;
      11'b01111000000 : romData <= 32'h0D000000;
      11'b01111000001 : romData <= 32'hF409639C;
      11'b01111000010 : romData <= 32'hADDE201A;
      11'b01111000011 : romData <= 32'hEFBE31AA;
      11'b01111000100 : romData <= 32'h00F08018;
      11'b01111000101 : romData <= 32'h00F06018;
      11'b01111000110 : romData <= 32'h00007086;
      11'b01111000111 : romData <= 32'h008813E4;
      11'b01111001000 : romData <= 32'h8C08849C;
      11'b01111001001 : romData <= 32'h08000010;
      11'b01111001010 : romData <= 32'hF409639C;
      11'b01111001011 : romData <= 32'h00F0A018;
      11'b01111001100 : romData <= 32'hAA19A59C;
      11'b01111001101 : romData <= 32'hD2FDFF07;
      11'b01111001110 : romData <= 32'h270040AB;
      11'b01111001111 : romData <= 32'h4AFFFF03;
      11'b01111010000 : romData <= 32'h00000015;
      11'b01111010001 : romData <= 32'h00F0A018;
      11'b01111010010 : romData <= 32'hC519A59C;
      11'b01111010011 : romData <= 32'hCCFDFF07;
      11'b01111010100 : romData <= 32'h00000015;
      11'b01111010101 : romData <= 32'h30000074;
      11'b01111010110 : romData <= 32'h43FFFF03;
      11'b01111010111 : romData <= 32'h270040AB;
      11'b01111011000 : romData <= 32'h5AFEFF07;
      11'b01111011001 : romData <= 32'h00000015;
      11'b01111011010 : romData <= 32'hFF006BA5;
      11'b01111011011 : romData <= 32'h6D0020AA;
      11'b01111011100 : romData <= 32'h00880BE4;
      11'b01111011101 : romData <= 32'h44010010;
      11'b01111011110 : romData <= 32'h00884BE4;
      11'b01111011111 : romData <= 32'h4E000010;
      11'b01111100000 : romData <= 32'h730020AA;
      11'b01111100001 : romData <= 32'h660020AA;
      11'b01111100010 : romData <= 32'h00880BE4;
      11'b01111100011 : romData <= 32'hE7000010;
      11'b01111100100 : romData <= 32'h00884BE4;
      11'b01111100101 : romData <= 32'h32000010;
      11'b01111100110 : romData <= 32'h680020AA;
      11'b01111100111 : romData <= 32'h630020AA;
      11'b01111101000 : romData <= 32'h00880BE4;
      11'b01111101001 : romData <= 32'hA6000010;
      11'b01111101010 : romData <= 32'h650020AA;
      11'b01111101011 : romData <= 32'h00880BE4;
      11'b01111101100 : romData <= 32'h2CFFFF0F;
      11'b01111101101 : romData <= 32'h00F0401B;
      11'b01111101110 : romData <= 32'h00F0001B;
      11'b01111101111 : romData <= 32'h8C085A9F;
      11'b01111110000 : romData <= 32'hF409189F;
      11'b01111110001 : romData <= 32'h00F0A018;
      11'b01111110010 : romData <= 32'h901BA59C;
      11'b01111110011 : romData <= 32'h04D09AE0;
      11'b01111110100 : romData <= 32'hABFDFF07;
      11'b01111110101 : romData <= 32'h04C078E0;
      11'b01111110110 : romData <= 32'h00F04018;
      11'b01111110111 : romData <= 32'h241BA29C;
      11'b01111111000 : romData <= 32'h0004201A;
      11'b01111111001 : romData <= 32'hFFFFE0AE;
      11'b01111111010 : romData <= 32'h00FC201B;
      11'b01111111011 : romData <= 32'h00054018;
      11'b01111111100 : romData <= 32'h00007186;
      11'b01111111101 : romData <= 32'h00B813E4;
      11'b01111111110 : romData <= 32'h12000010;
      11'b01111111111 : romData <= 32'h00C871E2;
      11'b10000000000 : romData <= 32'h009801D4;
      11'b10000000001 : romData <= 32'h04D09AE0;
      11'b10000000010 : romData <= 32'h04C078E0;
      11'b10000000011 : romData <= 32'h20B801D4;
      11'b10000000100 : romData <= 32'h1CC801D4;
      11'b10000000101 : romData <= 32'h188801D4;
      11'b10000000110 : romData <= 32'h0C2801D4;
      11'b10000000111 : romData <= 32'h98FDFF07;
      11'b10000001000 : romData <= 32'h149801D4;
      11'b10000001001 : romData <= 32'h14006186;
      11'b10000001010 : romData <= 32'h88FCFF07;
      11'b10000001011 : romData <= 32'h049873E0;
      11'b10000001100 : romData <= 32'h2000E186;
      11'b10000001101 : romData <= 32'h1C002187;
      11'b10000001110 : romData <= 32'h18002186;
      11'b10000001111 : romData <= 32'h0C00A184;
      11'b10000010000 : romData <= 32'h0400319E;
      11'b10000010001 : romData <= 32'h001031E4;
      11'b10000010010 : romData <= 32'hEAFFFF13;
      11'b10000010011 : romData <= 32'h00000015;
      11'b10000010100 : romData <= 32'h00F0A018;
      11'b10000010101 : romData <= 32'hBE000000;
      11'b10000010110 : romData <= 32'hAE1BA59C;
      11'b10000010111 : romData <= 32'h00880BE4;
      11'b10000011000 : romData <= 32'h44000010;
      11'b10000011001 : romData <= 32'h690020AA;
      11'b10000011010 : romData <= 32'h00880BE4;
      11'b10000011011 : romData <= 32'hFDFEFF0F;
      11'b10000011100 : romData <= 32'hADDE201A;
      11'b10000011101 : romData <= 32'hEFBE31AA;
      11'b10000011110 : romData <= 32'h00007086;
      11'b10000011111 : romData <= 32'h00F08018;
      11'b10000100000 : romData <= 32'h008813E4;
      11'b10000100001 : romData <= 32'h00F06018;
      11'b10000100010 : romData <= 32'h04003086;
      11'b10000100011 : romData <= 32'h8C08849C;
      11'b10000100100 : romData <= 32'h4F000010;
      11'b10000100101 : romData <= 32'hF409639C;
      11'b10000100110 : romData <= 32'h00F0A018;
      11'b10000100111 : romData <= 32'h048801D4;
      11'b10000101000 : romData <= 32'h000001D4;
      11'b10000101001 : romData <= 32'h76FDFF07;
      11'b10000101010 : romData <= 32'h0B1AA59C;
      11'b10000101011 : romData <= 32'hEEFEFF03;
      11'b10000101100 : romData <= 32'h270040AB;
      11'b10000101101 : romData <= 32'h00880BE4;
      11'b10000101110 : romData <= 32'h38000010;
      11'b10000101111 : romData <= 32'h00884BE4;
      11'b10000110000 : romData <= 32'h1E000010;
      11'b10000110001 : romData <= 32'h740020AA;
      11'b10000110010 : romData <= 32'h700020AA;
      11'b10000110011 : romData <= 32'h00880BE4;
      11'b10000110100 : romData <= 32'h36000010;
      11'b10000110101 : romData <= 32'h720020AA;
      11'b10000110110 : romData <= 32'h00880BE4;
      11'b10000110111 : romData <= 32'hE1FEFF0F;
      11'b10000111000 : romData <= 32'hADDE201A;
      11'b10000111001 : romData <= 32'h0004A01A;
      11'b10000111010 : romData <= 32'hEFBE31AA;
      11'b10000111011 : romData <= 32'h00007586;
      11'b10000111100 : romData <= 32'h008833E4;
      11'b10000111101 : romData <= 32'hE2000010;
      11'b10000111110 : romData <= 32'h00F0A018;
      11'b10000111111 : romData <= 32'h040035AA;
      11'b10001000000 : romData <= 32'h00007186;
      11'b10001000001 : romData <= 32'h020020AA;
      11'b10001000010 : romData <= 32'h088873E2;
      11'b10001000011 : romData <= 32'h0000201A;
      11'b10001000100 : romData <= 32'h009831E4;
      11'b10001000101 : romData <= 32'hD5000010;
      11'b10001000110 : romData <= 32'h0088F5E2;
      11'b10001000111 : romData <= 32'h00F0A018;
      11'b10001001000 : romData <= 32'h00F08018;
      11'b10001001001 : romData <= 32'h00F06018;
      11'b10001001010 : romData <= 32'h4C19A59C;
      11'b10001001011 : romData <= 32'h8C08849C;
      11'b10001001100 : romData <= 32'h87FFFF03;
      11'b10001001101 : romData <= 32'hF409639C;
      11'b10001001110 : romData <= 32'h00880BE4;
      11'b10001001111 : romData <= 32'h2D000010;
      11'b10001010000 : romData <= 32'h760020AA;
      11'b10001010001 : romData <= 32'h00880BE4;
      11'b10001010010 : romData <= 32'hC6FEFF0F;
      11'b10001010011 : romData <= 32'h00F0A018;
      11'b10001010100 : romData <= 32'h00F08018;
      11'b10001010101 : romData <= 32'h00F06018;
      11'b10001010110 : romData <= 32'hF619A59C;
      11'b10001010111 : romData <= 32'h8C08849C;
      11'b10001011000 : romData <= 32'h47FDFF07;
      11'b10001011001 : romData <= 32'hF409639C;
      11'b10001011010 : romData <= 32'hBEFEFF03;
      11'b10001011011 : romData <= 32'h0000C01B;
      11'b10001011100 : romData <= 32'h00F0A018;
      11'b10001011101 : romData <= 32'h00F06018;
      11'b10001011110 : romData <= 32'hC61BA59C;
      11'b10001011111 : romData <= 32'h00008018;
      11'b10001100000 : romData <= 32'h3FFDFF07;
      11'b10001100001 : romData <= 32'h8C08639C;
      11'b10001100010 : romData <= 32'h2CFEFF07;
      11'b10001100011 : romData <= 32'h270040AB;
      11'b10001100100 : romData <= 32'hB5FEFF03;
      11'b10001100101 : romData <= 32'h00000015;
      11'b10001100110 : romData <= 32'h61FCFF07;
      11'b10001100111 : romData <= 32'h270040AB;
      11'b10001101000 : romData <= 32'hB1FEFF03;
      11'b10001101001 : romData <= 32'h00000015;
      11'b10001101010 : romData <= 32'h00F0A018;
      11'b10001101011 : romData <= 32'h00F08018;
      11'b10001101100 : romData <= 32'h00F06018;
      11'b10001101101 : romData <= 32'hE219A59C;
      11'b10001101110 : romData <= 32'h8C08849C;
      11'b10001101111 : romData <= 32'h30FDFF07;
      11'b10001110000 : romData <= 32'hF409639C;
      11'b10001110001 : romData <= 32'hA7FEFF03;
      11'b10001110010 : romData <= 32'h0100C0AB;
      11'b10001110011 : romData <= 32'h020060AA;
      11'b10001110100 : romData <= 32'h089831E2;
      11'b10001110101 : romData <= 32'hFFFF319E;
      11'b10001110110 : romData <= 32'h00F0A018;
      11'b10001110111 : romData <= 32'h008801D4;
      11'b10001111000 : romData <= 32'h27FDFF07;
      11'b10001111001 : romData <= 32'h1F1AA59C;
      11'b10001111010 : romData <= 32'h9FFEFF03;
      11'b10001111011 : romData <= 32'h270040AB;
      11'b10001111100 : romData <= 32'h0000201A;
      11'b10001111101 : romData <= 32'h00F08018;
      11'b10001111110 : romData <= 32'h00F06018;
      11'b10001111111 : romData <= 32'h008830E4;
      11'b10010000000 : romData <= 32'h8C08849C;
      11'b10010000001 : romData <= 32'h08000010;
      11'b10010000010 : romData <= 32'hF409639C;
      11'b10010000011 : romData <= 32'h00F0A018;
      11'b10010000100 : romData <= 32'h1BFDFF07;
      11'b10010000101 : romData <= 32'h481AA59C;
      11'b10010000110 : romData <= 32'h0000C019;
      11'b10010000111 : romData <= 32'h91FEFF03;
      11'b10010001000 : romData <= 32'h0004001A;
      11'b10010001001 : romData <= 32'h00F0A018;
      11'b10010001010 : romData <= 32'h15FDFF07;
      11'b10010001011 : romData <= 32'h5B1AA59C;
      11'b10010001100 : romData <= 32'h0000C019;
      11'b10010001101 : romData <= 32'h8BFEFF03;
      11'b10010001110 : romData <= 32'h0000001A;
      11'b10010001111 : romData <= 32'h0000201A;
      11'b10010010000 : romData <= 32'h008810E4;
      11'b10010010001 : romData <= 32'h05000010;
      11'b10010010010 : romData <= 32'hADDE201A;
      11'b10010010011 : romData <= 32'h00F0A018;
      11'b10010010100 : romData <= 32'h29FFFF03;
      11'b10010010101 : romData <= 32'h6E1AA59C;
      11'b10010010110 : romData <= 32'hEFBE31AA;
      11'b10010010111 : romData <= 32'h00007086;
      11'b10010011000 : romData <= 32'h008813E4;
      11'b10010011001 : romData <= 32'h05000010;
      11'b10010011010 : romData <= 32'h3F00201A;
      11'b10010011011 : romData <= 32'h00F0A018;
      11'b10010011100 : romData <= 32'h21FFFF03;
      11'b10010011101 : romData <= 32'h901AA59C;
      11'b10010011110 : romData <= 32'hFFFF31AA;
      11'b10010011111 : romData <= 32'h04007086;
      11'b10010100000 : romData <= 32'h0088B3E4;
      11'b10010100001 : romData <= 32'h21000010;
      11'b10010100010 : romData <= 32'h00F0A018;
      11'b10010100011 : romData <= 32'h1AFFFF03;
      11'b10010100100 : romData <= 32'hAD1AA59C;
      11'b10010100101 : romData <= 32'h0088B8E2;
      11'b10010100110 : romData <= 32'h00007587;
      11'b10010100111 : romData <= 32'h00003887;
      11'b10010101000 : romData <= 32'h00C81BE4;
      11'b10010101001 : romData <= 32'h10000010;
      11'b10010101010 : romData <= 32'h048838E2;
      11'b10010101011 : romData <= 32'h00F06018;
      11'b10010101100 : romData <= 32'h0000B586;
      11'b10010101101 : romData <= 32'h04D0BAE0;
      11'b10010101110 : romData <= 32'h00003887;
      11'b10010101111 : romData <= 32'h041082E0;
      11'b10010110000 : romData <= 32'h08C801D4;
      11'b10010110001 : romData <= 32'h04A801D4;
      11'b10010110010 : romData <= 32'h008801D4;
      11'b10010110011 : romData <= 32'hF409639C;
      11'b10010110100 : romData <= 32'h14B801D4;
      11'b10010110101 : romData <= 32'hEAFCFF07;
      11'b10010110110 : romData <= 32'h0C9801D4;
      11'b10010110111 : romData <= 32'h1400E186;
      11'b10010111000 : romData <= 32'h0C006186;
      11'b10010111001 : romData <= 32'h0100739E;
      11'b10010111010 : romData <= 32'h0400189F;
      11'b10010111011 : romData <= 32'h00003786;
      11'b10010111100 : romData <= 32'h009851E4;
      11'b10010111101 : romData <= 32'hE8FFFF13;
      11'b10010111110 : romData <= 32'h0004201A;
      11'b10010111111 : romData <= 32'h00F0A018;
      11'b10011000000 : romData <= 32'hFDFEFF03;
      11'b10011000001 : romData <= 32'hF31AA59C;
      11'b10011000010 : romData <= 32'h00F0401B;
      11'b10011000011 : romData <= 32'h00F04018;
      11'b10011000100 : romData <= 32'h0000001B;
      11'b10011000101 : romData <= 32'h0000601A;
      11'b10011000110 : romData <= 32'h0400E0AA;
      11'b10011000111 : romData <= 32'hCD1A5A9F;
      11'b10011001000 : romData <= 32'hF3FFFF03;
      11'b10011001001 : romData <= 32'h8C08429C;
      11'b10011001010 : romData <= 32'h0000201A;
      11'b10011001011 : romData <= 32'h00F0401B;
      11'b10011001100 : romData <= 32'h00F0001B;
      11'b10011001101 : romData <= 32'h008810E4;
      11'b10011001110 : romData <= 32'h8C085A9F;
      11'b10011001111 : romData <= 32'h07000010;
      11'b10011010000 : romData <= 32'hF409189F;
      11'b10011010001 : romData <= 32'h00F0A018;
      11'b10011010010 : romData <= 32'h6E1AA59C;
      11'b10011010011 : romData <= 32'h04D09AE0;
      11'b10011010100 : romData <= 32'hF9FEFF03;
      11'b10011010101 : romData <= 32'h04C078E0;
      11'b10011010110 : romData <= 32'hADDE201A;
      11'b10011010111 : romData <= 32'hEFBE31AA;
      11'b10011011000 : romData <= 32'h00007086;
      11'b10011011001 : romData <= 32'h008813E4;
      11'b10011011010 : romData <= 32'h05000010;
      11'b10011011011 : romData <= 32'h3F00201A;
      11'b10011011100 : romData <= 32'h00F0A018;
      11'b10011011101 : romData <= 32'hF6FFFF03;
      11'b10011011110 : romData <= 32'h901AA59C;
      11'b10011011111 : romData <= 32'hFFFF31AA;
      11'b10011100000 : romData <= 32'h04007086;
      11'b10011100001 : romData <= 32'h0088B3E4;
      11'b10011100010 : romData <= 32'h04000010;
      11'b10011100011 : romData <= 32'h00F0A018;
      11'b10011100100 : romData <= 32'hEFFFFF03;
      11'b10011100101 : romData <= 32'hAD1AA59C;
      11'b10011100110 : romData <= 32'h00F0A018;
      11'b10011100111 : romData <= 32'h011BA59C;
      11'b10011101000 : romData <= 32'h04D09AE0;
      11'b10011101001 : romData <= 32'hB6FCFF07;
      11'b10011101010 : romData <= 32'h04C078E0;
      11'b10011101011 : romData <= 32'h00F0A018;
      11'b10011101100 : romData <= 32'h0004201A;
      11'b10011101101 : romData <= 32'h0000601A;
      11'b10011101110 : romData <= 32'h040040A8;
      11'b10011101111 : romData <= 32'hFFFFE0AE;
      11'b10011110000 : romData <= 32'h00FC201B;
      11'b10011110001 : romData <= 32'h241BA59C;
      11'b10011110010 : romData <= 32'h0000A286;
      11'b10011110011 : romData <= 32'h009855E4;
      11'b10011110100 : romData <= 32'h0D000010;
      11'b10011110101 : romData <= 32'h04D09AE0;
      11'b10011110110 : romData <= 32'h00F0A018;
      11'b10011110111 : romData <= 32'h4B1BA59C;
      11'b10011111000 : romData <= 32'hA7FCFF07;
      11'b10011111001 : romData <= 32'h04C078E0;
      11'b10011111010 : romData <= 32'h00006018;
      11'b10011111011 : romData <= 32'h00008284;
      11'b10011111100 : romData <= 32'h9DFBFF07;
      11'b10011111101 : romData <= 32'h00000015;
      11'b10011111110 : romData <= 32'h00F0A018;
      11'b10011111111 : romData <= 32'hD4FFFF03;
      11'b10100000000 : romData <= 32'h641BA59C;
      11'b10100000001 : romData <= 32'h0000B186;
      11'b10100000010 : romData <= 32'h00B815E4;
      11'b10100000011 : romData <= 32'h14000010;
      11'b10100000100 : romData <= 32'h00C8B1E2;
      11'b10100000101 : romData <= 32'h00A801D4;
      11'b10100000110 : romData <= 32'h04D09AE0;
      11'b10100000111 : romData <= 32'h04C078E0;
      11'b10100001000 : romData <= 32'h24B801D4;
      11'b10100001001 : romData <= 32'h209801D4;
      11'b10100001010 : romData <= 32'h1CC801D4;
      11'b10100001011 : romData <= 32'h188801D4;
      11'b10100001100 : romData <= 32'h0C2801D4;
      11'b10100001101 : romData <= 32'h92FCFF07;
      11'b10100001110 : romData <= 32'h14A801D4;
      11'b10100001111 : romData <= 32'h1400A186;
      11'b10100010000 : romData <= 32'h82FBFF07;
      11'b10100010001 : romData <= 32'h04A875E0;
      11'b10100010010 : romData <= 32'h2400E186;
      11'b10100010011 : romData <= 32'h20006186;
      11'b10100010100 : romData <= 32'h1C002187;
      11'b10100010101 : romData <= 32'h18002186;
      11'b10100010110 : romData <= 32'h0C00A184;
      11'b10100010111 : romData <= 32'h0100739E;
      11'b10100011000 : romData <= 32'hDAFFFF03;
      11'b10100011001 : romData <= 32'h0400319E;
      11'b10100011010 : romData <= 32'h0000F786;
      11'b10100011011 : romData <= 32'h0400319E;
      11'b10100011100 : romData <= 32'hFCBFF1D7;
      11'b10100011101 : romData <= 32'h28FFFF03;
      11'b10100011110 : romData <= 32'h009831E4;
      11'b10100011111 : romData <= 32'h9EFEFF03;
      11'b10100100000 : romData <= 32'h7A1BA59C;
      11'b10100100001 : romData <= 32'h00F0401B;
      11'b10100100010 : romData <= 32'h00F0001B;
      11'b10100100011 : romData <= 32'h8C085A9F;
      11'b10100100100 : romData <= 32'hF409189F;
      11'b10100100101 : romData <= 32'h00F0A018;
      11'b10100100110 : romData <= 32'hC91BA59C;
      11'b10100100111 : romData <= 32'h04D09AE0;
      11'b10100101000 : romData <= 32'h77FCFF07;
      11'b10100101001 : romData <= 32'h04C078E0;
      11'b10100101010 : romData <= 32'h00F0C019;
      11'b10100101011 : romData <= 32'hEB1B2E9E;
      11'b10100101100 : romData <= 32'h00004018;
      11'b10100101101 : romData <= 32'h0C8801D4;
      11'b10100101110 : romData <= 32'h04D09AE0;
      11'b10100101111 : romData <= 32'h04C078E0;
      11'b10100110000 : romData <= 32'h6FFCFF07;
      11'b10100110001 : romData <= 32'h0C00A184;
      11'b10100110010 : romData <= 32'h0000201A;
      11'b10100110011 : romData <= 32'h0002601A;
      11'b10100110100 : romData <= 32'h0200A0AA;
      11'b10100110101 : romData <= 32'h00A802E4;
      11'b10100110110 : romData <= 32'h03000010;
      11'b10100110111 : romData <= 32'h00000015;
      11'b10100111000 : romData <= 32'h0100F172;
      11'b10100111001 : romData <= 32'h008811D4;
      11'b10100111010 : romData <= 32'h0400319E;
      11'b10100111011 : romData <= 32'h009831E4;
      11'b10100111100 : romData <= 32'hF9FFFF13;
      11'b10100111101 : romData <= 32'h0200A0AA;
      11'b10100111110 : romData <= 32'h00F0A018;
      11'b10100111111 : romData <= 32'hF71BA59C;
      11'b10101000000 : romData <= 32'h04D09AE0;
      11'b10101000001 : romData <= 32'h5EFCFF07;
      11'b10101000010 : romData <= 32'h04C078E0;
      11'b10101000011 : romData <= 32'h0000201A;
      11'b10101000100 : romData <= 32'h0000C019;
      11'b10101000101 : romData <= 32'h1D0020AB;
      11'b10101000110 : romData <= 32'h0002E01A;
      11'b10101000111 : romData <= 32'h020060AA;
      11'b10101001000 : romData <= 32'h009802E4;
      11'b10101001001 : romData <= 32'h03000010;
      11'b10101001010 : romData <= 32'h00000015;
      11'b10101001011 : romData <= 32'h01007173;
      11'b10101001100 : romData <= 32'h00007187;
      11'b10101001101 : romData <= 32'h00881BE4;
      11'b10101001110 : romData <= 32'h13000010;
      11'b10101001111 : romData <= 32'h00C84EE4;
      11'b10101010000 : romData <= 32'h10000010;
      11'b10101010001 : romData <= 32'h00000015;
      11'b10101010010 : romData <= 32'h00007187;
      11'b10101010011 : romData <= 32'h04D09AE0;
      11'b10101010100 : romData <= 32'h088801D4;
      11'b10101010101 : romData <= 32'h008801D4;
      11'b10101010110 : romData <= 32'h04D801D4;
      11'b10101010111 : romData <= 32'h04C078E0;
      11'b10101011000 : romData <= 32'h1CC801D4;
      11'b10101011001 : romData <= 32'h18B801D4;
      11'b10101011010 : romData <= 32'h148801D4;
      11'b10101011011 : romData <= 32'h44FCFF07;
      11'b10101011100 : romData <= 32'h1000A184;
      11'b10101011101 : romData <= 32'h1C002187;
      11'b10101011110 : romData <= 32'h1800E186;
      11'b10101011111 : romData <= 32'h14002186;
      11'b10101100000 : romData <= 32'h0100CE9D;
      11'b10101100001 : romData <= 32'h0400319E;
      11'b10101100010 : romData <= 32'h00B831E4;
      11'b10101100011 : romData <= 32'hE5FFFF13;
      11'b10101100100 : romData <= 32'h020060AA;
      11'b10101100101 : romData <= 32'h0000201A;
      11'b10101100110 : romData <= 32'h00880EE4;
      11'b10101100111 : romData <= 32'h10000010;
      11'b10101101000 : romData <= 32'h030020AA;
      11'b10101101001 : romData <= 32'h00F0A018;
      11'b10101101010 : romData <= 32'h007001D4;
      11'b10101101011 : romData <= 32'h211CA59C;
      11'b10101101100 : romData <= 32'h04D09AE0;
      11'b10101101101 : romData <= 32'h32FCFF07;
      11'b10101101110 : romData <= 32'h04C078E0;
      11'b10101101111 : romData <= 32'h00F0A018;
      11'b10101110000 : romData <= 32'h007001D4;
      11'b10101110001 : romData <= 32'h3A1CA59C;
      11'b10101110010 : romData <= 32'h04D09AE0;
      11'b10101110011 : romData <= 32'h2CFCFF07;
      11'b10101110100 : romData <= 32'h04C078E0;
      11'b10101110101 : romData <= 32'hA3FDFF03;
      11'b10101110110 : romData <= 32'h0000C019;
      11'b10101110111 : romData <= 32'h0100429C;
      11'b10101111000 : romData <= 32'h008822E4;
      11'b10101111001 : romData <= 32'hB6FFFF13;
      11'b10101111010 : romData <= 32'h04D09AE0;
      11'b10101111011 : romData <= 32'hF5FFFF03;
      11'b10101111100 : romData <= 32'h00F0A018;
      11'b10101111101 : romData <= 32'hB5FCFF07;
      11'b10101111110 : romData <= 32'h270040AB;
      11'b10101111111 : romData <= 32'hB3FCFF07;
      11'b10110000000 : romData <= 32'hFF000BA7;
      11'b10110000001 : romData <= 32'hD0FF189F;
      11'b10110000010 : romData <= 32'h020020AA;
      11'b10110000011 : romData <= 32'h088838E2;
      11'b10110000100 : romData <= 32'hFF004BA6;
      11'b10110000101 : romData <= 32'h00C031E2;
      11'b10110000110 : romData <= 32'h008831E2;
      11'b10110000111 : romData <= 32'hD0FF529E;
      11'b10110001000 : romData <= 32'h91FDFF03;
      11'b10110001001 : romData <= 32'h008852E2;
      11'b10110001010 : romData <= 32'h551CA59C;
      11'b10110001011 : romData <= 32'h34FEFF03;
      11'b10110001100 : romData <= 32'h00008018;
      11'b10110001101 : romData <= 32'h18000010;
      11'b10110001110 : romData <= 32'h080020AA;
      11'b10110001111 : romData <= 32'h0888D6E2;
      11'b10110010000 : romData <= 32'h01009C9F;
      11'b10110010001 : romData <= 32'h040020AA;
      11'b10110010010 : romData <= 32'h00883CE4;
      11'b10110010011 : romData <= 32'h30000010;
      11'b10110010100 : romData <= 32'h00B0C2E2;
      11'b10110010101 : romData <= 32'h0000201A;
      11'b10110010110 : romData <= 32'h008810E4;
      11'b10110010111 : romData <= 32'h10000010;
      11'b10110011000 : romData <= 32'h0000601A;
      11'b10110011001 : romData <= 32'h008834E4;
      11'b10110011010 : romData <= 32'h7EFDFF13;
      11'b10110011011 : romData <= 32'h010040AA;
      11'b10110011100 : romData <= 32'h00F0A018;
      11'b10110011101 : romData <= 32'h00F08018;
      11'b10110011110 : romData <= 32'h00F06018;
      11'b10110011111 : romData <= 32'h631CA59C;
      11'b10110100000 : romData <= 32'h8C08849C;
      11'b10110100001 : romData <= 32'hFEFBFF07;
      11'b10110100010 : romData <= 32'hF409639C;
      11'b10110100011 : romData <= 32'h75FDFF03;
      11'b10110100100 : romData <= 32'h049092E2;
      11'b10110100101 : romData <= 32'hEBFFFF03;
      11'b10110100110 : romData <= 32'h0000C01A;
      11'b10110100111 : romData <= 32'h020020AA;
      11'b10110101000 : romData <= 32'h088894E3;
      11'b10110101001 : romData <= 32'hFF3F34A6;
      11'b10110101010 : romData <= 32'h009831E4;
      11'b10110101011 : romData <= 32'h07000010;
      11'b10110101100 : romData <= 32'h00F0A018;
      11'b10110101101 : romData <= 32'h00E001D4;
      11'b10110101110 : romData <= 32'h841CA59C;
      11'b10110101111 : romData <= 32'h00008018;
      11'b10110110000 : romData <= 32'hEFFBFF07;
      11'b10110110001 : romData <= 32'h04C078E0;
      11'b10110110010 : romData <= 32'h0000201A;
      11'b10110110011 : romData <= 32'h00881EE4;
      11'b10110110100 : romData <= 32'h11000010;
      11'b10110110101 : romData <= 32'h00E030E2;
      11'b10110110110 : romData <= 32'h01007672;
      11'b10110110111 : romData <= 32'h009811D4;
      11'b10110111000 : romData <= 32'h0100949E;
      11'b10110111001 : romData <= 32'h00A06EE4;
      11'b10110111010 : romData <= 32'h09000010;
      11'b10110111011 : romData <= 32'h0000801B;
      11'b10110111100 : romData <= 32'h0000201A;
      11'b10110111101 : romData <= 32'h00881EE4;
      11'b10110111110 : romData <= 32'h05000010;
      11'b10110111111 : romData <= 32'h00000015;
      11'b10111000000 : romData <= 32'h04A010D4;
      11'b10111000001 : romData <= 32'h04A0D4E1;
      11'b10111000010 : romData <= 32'h0000801B;
      11'b10111000011 : romData <= 32'hD8FDFF03;
      11'b10111000100 : romData <= 32'hFFFF529E;
      11'b10111000101 : romData <= 32'h00003186;
      11'b10111000110 : romData <= 32'h01003172;
      11'b10111000111 : romData <= 32'h008816E4;
      11'b10111001000 : romData <= 32'hF0FFFF13;
      11'b10111001001 : romData <= 32'h04D0BAE0;
      11'b10111001010 : romData <= 32'h08B001D4;
      11'b10111001011 : romData <= 32'h048801D4;
      11'b10111001100 : romData <= 32'h00E001D4;
      11'b10111001101 : romData <= 32'h00008018;
      11'b10111001110 : romData <= 32'hD1FBFF07;
      11'b10111001111 : romData <= 32'h04C078E0;
      11'b10111010000 : romData <= 32'hE9FFFF03;
      11'b10111010001 : romData <= 32'h0100949E;
      11'b10111010010 : romData <= 32'h000004E4;
      11'b10111010011 : romData <= 32'h000060A9;
      11'b10111010100 : romData <= 32'h15000010;
      11'b10111010101 : romData <= 32'h000083A9;
      11'b10111010110 : romData <= 32'h0100C0A8;
      11'b10111010111 : romData <= 32'h000084E5;
      11'b10111011000 : romData <= 32'h05000010;
      11'b10111011001 : romData <= 32'h006084E4;
      11'b10111011010 : romData <= 32'h002084E0;
      11'b10111011011 : romData <= 32'hFCFFFF13;
      11'b10111011100 : romData <= 32'h0030C6E0;
      11'b10111011101 : romData <= 32'h0030EBE0;
      11'b10111011110 : romData <= 32'h4100C6B8;
      11'b10111011111 : romData <= 32'h02200CE1;
      11'b10111100000 : romData <= 32'h0060A4E4;
      11'b10111100001 : romData <= 32'h410084B8;
      11'b10111100010 : romData <= 32'h0400000C;
      11'b10111100011 : romData <= 32'h00000015;
      11'b10111100100 : romData <= 32'h000067A9;
      11'b10111100101 : romData <= 32'h000088A9;
      11'b10111100110 : romData <= 32'h000026E4;
      11'b10111100111 : romData <= 32'hF7FFFF13;
      11'b10111101000 : romData <= 32'h0030EBE0;
      11'b10111101001 : romData <= 32'h00480044;
      11'b10111101010 : romData <= 32'h00000015;
      11'b10111101011 : romData <= 32'h0000A9A9;
      11'b10111101100 : romData <= 32'hE6FFFF07;
      11'b10111101101 : romData <= 32'h00000015;
      11'b10111101110 : romData <= 32'h00680044;
      11'b10111101111 : romData <= 32'h00006CA9;
      11'b10111110000 : romData <= 32'h65202449;
      11'b10111110001 : romData <= 32'h726F7272;
      11'b10111110010 : romData <= 32'h44000A21;
      11'b10111110011 : romData <= 32'h72652024;
      11'b10111110100 : romData <= 32'h0A726F72;
      11'b10111110101 : romData <= 32'h71726900;
      11'b10111110110 : romData <= 32'h3F3F000A;
      11'b10111110111 : romData <= 32'h73000A3F;
      11'b10111111000 : romData <= 32'h65747379;
      11'b10111111001 : romData <= 32'h000A216D;
      11'b10111111010 : romData <= 32'h63656843;
      11'b10111111011 : romData <= 32'h676E696B;
      11'b10111111100 : romData <= 32'h73616C20;
      11'b10111111101 : romData <= 32'h61702074;
      11'b10111111110 : romData <= 32'h6F206567;
      11'b10111111111 : romData <= 32'h6C662066;
      11'b11000000000 : romData <= 32'h20687361;
      11'b11000000001 : romData <= 32'h74706D65;
      11'b11000000010 : romData <= 32'h46000A79;
      11'b11000000011 : romData <= 32'h6873616C;
      11'b11000000100 : romData <= 32'h72726520;
      11'b11000000101 : romData <= 32'h0A21726F;
      11'b11000000110 : romData <= 32'h61724500;
      11'b11000000111 : romData <= 32'h676E6973;
      11'b11000001000 : romData <= 32'h73616C20;
      11'b11000001001 : romData <= 32'h61702074;
      11'b11000001010 : romData <= 32'h6F206567;
      11'b11000001011 : romData <= 32'h6C462066;
      11'b11000001100 : romData <= 32'h0A687361;
      11'b11000001101 : romData <= 32'h69725700;
      11'b11000001110 : romData <= 32'h676E6974;
      11'b11000001111 : romData <= 32'h73657420;
      11'b11000010000 : romData <= 32'h65732074;
      11'b11000010001 : romData <= 32'h6E657571;
      11'b11000010010 : romData <= 32'h74206563;
      11'b11000010011 : romData <= 32'h6C66206F;
      11'b11000010100 : romData <= 32'h2E687361;
      11'b11000010101 : romData <= 32'h6556000A;
      11'b11000010110 : romData <= 32'h79666972;
      11'b11000010111 : romData <= 32'h20676E69;
      11'b11000011000 : romData <= 32'h74736574;
      11'b11000011001 : romData <= 32'h71657320;
      11'b11000011010 : romData <= 32'h636E6575;
      11'b11000011011 : romData <= 32'h72662065;
      11'b11000011100 : romData <= 32'h66206D6F;
      11'b11000011101 : romData <= 32'h6873616C;
      11'b11000011110 : romData <= 32'h54000A2E;
      11'b11000011111 : romData <= 32'h20747365;
      11'b11000100000 : romData <= 32'h6C696166;
      11'b11000100001 : romData <= 32'h203A6465;
      11'b11000100010 : romData <= 32'h3A206425;
      11'b11000100011 : romData <= 32'h25783020;
      11'b11000100100 : romData <= 32'h3D2F2058;
      11'b11000100101 : romData <= 32'h25783020;
      11'b11000100110 : romData <= 32'h46000A58;
      11'b11000100111 : romData <= 32'h6873616C;
      11'b11000101000 : romData <= 32'h73657420;
      11'b11000101001 : romData <= 32'h6B6F2074;
      11'b11000101010 : romData <= 32'h0A2E7961;
      11'b11000101011 : romData <= 32'h5343000A;
      11'b11000101100 : romData <= 32'h3637342D;
      11'b11000101101 : romData <= 32'h626D4520;
      11'b11000101110 : romData <= 32'h65646465;
      11'b11000101111 : romData <= 32'h79532064;
      11'b11000110000 : romData <= 32'h6D657473;
      11'b11000110001 : romData <= 32'h73654420;
      11'b11000110010 : romData <= 32'h0A6E6769;
      11'b11000110011 : romData <= 32'h65704F00;
      11'b11000110100 : romData <= 32'h7369726E;
      11'b11000110101 : romData <= 32'h61622063;
      11'b11000110110 : romData <= 32'h20646573;
      11'b11000110111 : romData <= 32'h74726976;
      11'b11000111000 : romData <= 32'h206C6175;
      11'b11000111001 : romData <= 32'h746F7250;
      11'b11000111010 : romData <= 32'h7079746F;
      11'b11000111011 : romData <= 32'h000A2E65;
      11'b11000111100 : romData <= 32'h6C697542;
      11'b11000111101 : romData <= 32'h65762064;
      11'b11000111110 : romData <= 32'h6F697372;
      11'b11000111111 : romData <= 32'h44203A6E;
      11'b11001000000 : romData <= 32'h33312069;
      11'b11001000001 : romData <= 32'h62654620;
      11'b11001000010 : romData <= 32'h32303220;
      11'b11001000011 : romData <= 32'h30312034;
      11'b11001000100 : romData <= 32'h3A37323A;
      11'b11001000101 : romData <= 32'h43203235;
      11'b11001000110 : romData <= 32'h0A0A5445;
      11'b11001000111 : romData <= 32'h61204900;
      11'b11001001000 : romData <= 32'h5043206D;
      11'b11001001001 : romData <= 32'h64252055;
      11'b11001001010 : romData <= 32'h20666F20;
      11'b11001001011 : romData <= 32'h72206425;
      11'b11001001100 : romData <= 32'h696E6E75;
      11'b11001001101 : romData <= 32'h6120676E;
      11'b11001001110 : romData <= 32'h25002074;
      11'b11001001111 : romData <= 32'h2E642564;
      11'b11001010000 : romData <= 32'h64256425;
      11'b11001010001 : romData <= 32'h7A484D20;
      11'b11001010010 : romData <= 32'h000A0A2E;
      11'b11001010011 : romData <= 32'h63657845;
      11'b11001010100 : romData <= 32'h6E697475;
      11'b11001010101 : romData <= 32'h6C662067;
      11'b11001010110 : romData <= 32'h20687361;
      11'b11001010111 : romData <= 32'h676F7270;
      11'b11001011000 : romData <= 32'h2E6D6172;
      11'b11001011001 : romData <= 32'h000A2E2E;
      11'b11001011010 : romData <= 32'h6E776F44;
      11'b11001011011 : romData <= 32'h64616F6C;
      11'b11001011100 : romData <= 32'h6F64203A;
      11'b11001011101 : romData <= 32'h000A656E;
      11'b11001011110 : romData <= 32'h64616552;
      11'b11001011111 : romData <= 32'h20676E69;
      11'b11001100000 : romData <= 32'h65646F63;
      11'b11001100001 : romData <= 32'h62617420;
      11'b11001100010 : romData <= 32'h000A656C;
      11'b11001100011 : romData <= 32'h6E776F44;
      11'b11001100100 : romData <= 32'h64616F6C;
      11'b11001100101 : romData <= 32'h6573203A;
      11'b11001100110 : romData <= 32'h64612074;
      11'b11001100111 : romData <= 32'h73657264;
      11'b11001101000 : romData <= 32'h203D2073;
      11'b11001101001 : romData <= 32'h58257830;
      11'b11001101010 : romData <= 32'h7245000A;
      11'b11001101011 : romData <= 32'h2C726F72;
      11'b11001101100 : romData <= 32'h206F6E20;
      11'b11001101101 : romData <= 32'h676F7270;
      11'b11001101110 : romData <= 32'h206D6172;
      11'b11001101111 : romData <= 32'h64616F6C;
      11'b11001110000 : romData <= 32'h0A216465;
      11'b11001110001 : romData <= 32'h65784500;
      11'b11001110010 : romData <= 32'h69747563;
      11'b11001110011 : romData <= 32'h6C20676E;
      11'b11001110100 : romData <= 32'h6564616F;
      11'b11001110101 : romData <= 32'h72702064;
      11'b11001110110 : romData <= 32'h6172676F;
      11'b11001110111 : romData <= 32'h2E2E2E6D;
      11'b11001111000 : romData <= 32'h6553000A;
      11'b11001111001 : romData <= 32'h6E697474;
      11'b11001111010 : romData <= 32'h72702067;
      11'b11001111011 : romData <= 32'h202E676F;
      11'b11001111100 : romData <= 32'h65646F6D;
      11'b11001111101 : romData <= 32'h6553000A;
      11'b11001111110 : romData <= 32'h6E697474;
      11'b11001111111 : romData <= 32'h65762067;
      11'b11010000000 : romData <= 32'h2E666972;
      11'b11010000001 : romData <= 32'h646F6D20;
      11'b11010000010 : romData <= 32'h4E000A65;
      11'b11010000011 : romData <= 32'h7270206F;
      11'b11010000100 : romData <= 32'h6172676F;
      11'b11010000101 : romData <= 32'h7270206D;
      11'b11010000110 : romData <= 32'h6E657365;
      11'b11010000111 : romData <= 32'h50000A74;
      11'b11010001000 : romData <= 32'h72676F72;
      11'b11010001001 : romData <= 32'h69206D61;
      11'b11010001010 : romData <= 32'h656D206E;
      11'b11010001011 : romData <= 32'h7266206D;
      11'b11010001100 : romData <= 32'h62206D6F;
      11'b11010001101 : romData <= 32'h2B657361;
      11'b11010001110 : romData <= 32'h6F742030;
      11'b11010001111 : romData <= 32'h73616220;
      11'b11010010000 : romData <= 32'h78302B65;
      11'b11010010001 : romData <= 32'h000A5825;
      11'b11010010010 : romData <= 32'h74697753;
      11'b11010010011 : romData <= 32'h64656863;
      11'b11010010100 : romData <= 32'h206F7420;
      11'b11010010101 : romData <= 32'h73616C46;
      11'b11010010110 : romData <= 32'h53000A68;
      11'b11010010111 : romData <= 32'h63746977;
      11'b11010011000 : romData <= 32'h20646568;
      11'b11010011001 : romData <= 32'h53206F74;
      11'b11010011010 : romData <= 32'h6D615244;
      11'b11010011011 : romData <= 32'h6C50000A;
      11'b11010011100 : romData <= 32'h65736165;
      11'b11010011101 : romData <= 32'h61686320;
      11'b11010011110 : romData <= 32'h2065676E;
      11'b11010011111 : romData <= 32'h74206F74;
      11'b11010100000 : romData <= 32'h53206568;
      11'b11010100001 : romData <= 32'h4D415244;
      11'b11010100010 : romData <= 32'h20796220;
      11'b11010100011 : romData <= 32'h000A742A;
      11'b11010100100 : romData <= 32'h70206F4E;
      11'b11010100101 : romData <= 32'h72676F72;
      11'b11010100110 : romData <= 32'h6C206D61;
      11'b11010100111 : romData <= 32'h6564616F;
      11'b11010101000 : romData <= 32'h6E692064;
      11'b11010101001 : romData <= 32'h52445320;
      11'b11010101010 : romData <= 32'h0A216D61;
      11'b11010101011 : romData <= 32'h6F725000;
      11'b11010101100 : romData <= 32'h6D617267;
      11'b11010101101 : romData <= 32'h656F6420;
      11'b11010101110 : romData <= 32'h6F6E2073;
      11'b11010101111 : romData <= 32'h69662074;
      11'b11010110000 : romData <= 32'h6E692074;
      11'b11010110001 : romData <= 32'h616C4620;
      11'b11010110010 : romData <= 32'h0A216873;
      11'b11010110011 : romData <= 32'h6D6F4300;
      11'b11010110100 : romData <= 32'h65726170;
      11'b11010110101 : romData <= 32'h72726520;
      11'b11010110110 : romData <= 32'h6120726F;
      11'b11010110111 : romData <= 32'h78302074;
      11'b11010111000 : romData <= 32'h3A205825;
      11'b11010111001 : romData <= 32'h25783020;
      11'b11010111010 : romData <= 32'h3D212058;
      11'b11010111011 : romData <= 32'h25783020;
      11'b11010111100 : romData <= 32'h43000A58;
      11'b11010111101 : romData <= 32'h61706D6F;
      11'b11010111110 : romData <= 32'h64206572;
      11'b11010111111 : romData <= 32'h0A656E6F;
      11'b11011000000 : romData <= 32'h65684300;
      11'b11011000001 : romData <= 32'h6E696B63;
      11'b11011000010 : romData <= 32'h66692067;
      11'b11011000011 : romData <= 32'h65687420;
      11'b11011000100 : romData <= 32'h616C6620;
      11'b11011000101 : romData <= 32'h69206873;
      11'b11011000110 : romData <= 32'h6D652073;
      11'b11011000111 : romData <= 32'h2E797470;
      11'b11011001000 : romData <= 32'h000A2E2E;
      11'b11011001001 : romData <= 32'h72617453;
      11'b11011001010 : romData <= 32'h6C662074;
      11'b11011001011 : romData <= 32'h20687361;
      11'b11011001100 : romData <= 32'h73617265;
      11'b11011001101 : romData <= 32'h79632065;
      11'b11011001110 : romData <= 32'h20656C63;
      11'b11011001111 : romData <= 32'h20726F66;
      11'b11011010000 : romData <= 32'h65676170;
      11'b11011010001 : romData <= 32'h25783020;
      11'b11011010010 : romData <= 32'h53000A58;
      11'b11011010011 : romData <= 32'h74726174;
      11'b11011010100 : romData <= 32'h6F727020;
      11'b11011010101 : romData <= 32'h6D617267;
      11'b11011010110 : romData <= 32'h676E696D;
      11'b11011010111 : romData <= 32'h616C6620;
      11'b11011011000 : romData <= 32'h000A6873;
      11'b11011011001 : romData <= 32'h676F7250;
      11'b11011011010 : romData <= 32'h6D6D6172;
      11'b11011011011 : romData <= 32'h20676E69;
      11'b11011011100 : romData <= 32'h696E6966;
      11'b11011011101 : romData <= 32'h64656873;
      11'b11011011110 : romData <= 32'h6F4E000A;
      11'b11011011111 : romData <= 32'h6F727020;
      11'b11011100000 : romData <= 32'h6D617267;
      11'b11011100001 : romData <= 32'h206E6920;
      11'b11011100010 : romData <= 32'h73616C66;
      11'b11011100011 : romData <= 32'h000A2168;
      11'b11011100100 : romData <= 32'h63656843;
      11'b11011100101 : romData <= 32'h676E696B;
      11'b11011100110 : romData <= 32'h20666920;
      11'b11011100111 : romData <= 32'h73616C66;
      11'b11011101000 : romData <= 32'h73692068;
      11'b11011101001 : romData <= 32'h69642720;
      11'b11011101010 : romData <= 32'h27797472;
      11'b11011101011 : romData <= 32'h6C46000A;
      11'b11011101100 : romData <= 32'h20687361;
      11'b11011101101 : romData <= 32'h65207369;
      11'b11011101110 : romData <= 32'h7974706D;
      11'b11011101111 : romData <= 32'h72652820;
      11'b11011110000 : romData <= 32'h64657361;
      11'b11011110001 : romData <= 32'h0A0A2E29;
      11'b11011110010 : romData <= 32'h61745300;
      11'b11011110011 : romData <= 32'h6E697472;
      11'b11011110100 : romData <= 32'h69732067;
      11'b11011110101 : romData <= 32'h656C706D;
      11'b11011110110 : romData <= 32'h52445320;
      11'b11011110111 : romData <= 32'h6D206D61;
      11'b11011111000 : romData <= 32'h68636D65;
      11'b11011111001 : romData <= 32'h2E6B6365;
      11'b11011111010 : romData <= 32'h57000A0A;
      11'b11011111011 : romData <= 32'h69746972;
      11'b11011111100 : romData <= 32'h2E2E676E;
      11'b11011111101 : romData <= 32'h56000A2E;
      11'b11011111110 : romData <= 32'h66697265;
      11'b11011111111 : romData <= 32'h676E6979;
      11'b11100000000 : romData <= 32'h0A2E2E2E;
      11'b11100000001 : romData <= 32'h72724500;
      11'b11100000010 : romData <= 32'h4020726F;
      11'b11100000011 : romData <= 32'h58257830;
      11'b11100000100 : romData <= 32'h30203A20;
      11'b11100000101 : romData <= 32'h20582578;
      11'b11100000110 : romData <= 32'h30203D21;
      11'b11100000111 : romData <= 32'h0A582578;
      11'b11100001000 : romData <= 32'h20724E00;
      11'b11100001001 : romData <= 32'h6520666F;
      11'b11100001010 : romData <= 32'h726F7272;
      11'b11100001011 : romData <= 32'h6F662073;
      11'b11100001100 : romData <= 32'h20646E75;
      11'b11100001101 : romData <= 32'h6425203A;
      11'b11100001110 : romData <= 32'h654D000A;
      11'b11100001111 : romData <= 32'h6568636D;
      11'b11100010000 : romData <= 32'h64206B63;
      11'b11100010001 : romData <= 32'h2C656E6F;
      11'b11100010010 : romData <= 32'h20642520;
      11'b11100010011 : romData <= 32'h6F727265;
      11'b11100010100 : romData <= 32'h0A0A7372;
      11'b11100010101 : romData <= 32'h6B6E5500;
      11'b11100010110 : romData <= 32'h6E776F6E;
      11'b11100010111 : romData <= 32'h646F6320;
      11'b11100011000 : romData <= 32'h43002165;
      11'b11100011001 : romData <= 32'h6F6E6E61;
      11'b11100011010 : romData <= 32'h72702074;
      11'b11100011011 : romData <= 32'h6172676F;
      11'b11100011100 : romData <= 32'h6C66206D;
      11'b11100011101 : romData <= 32'h2C687361;
      11'b11100011110 : romData <= 32'h6F626120;
      11'b11100011111 : romData <= 32'h6E697472;
      11'b11100100000 : romData <= 32'h000A2167;
      11'b11100100001 : romData <= 32'h6E776F44;
      11'b11100100010 : romData <= 32'h64616F6C;
      11'b11100100011 : romData <= 32'h7461203A;
      11'b11100100100 : romData <= 32'h25783020;
      11'b11100100101 : romData <= 32'h56000A58;
      11'b11100100110 : romData <= 32'h66697265;
      11'b11100100111 : romData <= 32'h74616369;
      11'b11100101000 : romData <= 32'h206E6F69;
      11'b11100101001 : romData <= 32'h6F727265;
      11'b11100101010 : romData <= 32'h74612072;
      11'b11100101011 : romData <= 32'h25783020;
      11'b11100101100 : romData <= 32'h203A2058;
      11'b11100101101 : romData <= 32'h58257830;
      11'b11100101110 : romData <= 32'h203D2120;
      11'b11100101111 : romData <= 32'h58257830;
      11'b11100110000 : romData <= 32'h6E4B000A;
      11'b11100110001 : romData <= 32'h206E776F;
      11'b11100110010 : romData <= 32'h33325352;
      11'b11100110011 : romData <= 32'h6F632032;
      11'b11100110100 : romData <= 32'h6E616D6D;
      11'b11100110101 : romData <= 32'h0A3A7364;
      11'b11100110110 : romData <= 32'h20202400;
      11'b11100110111 : romData <= 32'h72617453;
      11'b11100111000 : romData <= 32'h68742074;
      11'b11100111001 : romData <= 32'h72702065;
      11'b11100111010 : romData <= 32'h6172676F;
      11'b11100111011 : romData <= 32'h6F6C206D;
      11'b11100111100 : romData <= 32'h64656461;
      11'b11100111101 : romData <= 32'h206E6920;
      11'b11100111110 : romData <= 32'h67726174;
      11'b11100111111 : romData <= 32'h000A7465;
      11'b11101000000 : romData <= 32'h5320702A;
      11'b11101000001 : romData <= 32'h70207465;
      11'b11101000010 : romData <= 32'h72676F72;
      11'b11101000011 : romData <= 32'h696D6D61;
      11'b11101000100 : romData <= 32'h6D20676E;
      11'b11101000101 : romData <= 32'h2065646F;
      11'b11101000110 : romData <= 32'h66656428;
      11'b11101000111 : romData <= 32'h746C7561;
      11'b11101001000 : romData <= 32'h2A000A29;
      11'b11101001001 : romData <= 32'h65532076;
      11'b11101001010 : romData <= 32'h65762074;
      11'b11101001011 : romData <= 32'h69666972;
      11'b11101001100 : romData <= 32'h69746163;
      11'b11101001101 : romData <= 32'h6D206E6F;
      11'b11101001110 : romData <= 32'h0A65646F;
      11'b11101001111 : romData <= 32'h20692A00;
      11'b11101010000 : romData <= 32'h776F6853;
      11'b11101010001 : romData <= 32'h666E6920;
      11'b11101010010 : romData <= 32'h6E6F206F;
      11'b11101010011 : romData <= 32'h6F727020;
      11'b11101010100 : romData <= 32'h6D617267;
      11'b11101010101 : romData <= 32'h206E6920;
      11'b11101010110 : romData <= 32'h67726174;
      11'b11101010111 : romData <= 32'h000A7465;
      11'b11101011000 : romData <= 32'h5420742A;
      11'b11101011001 : romData <= 32'h6C67676F;
      11'b11101011010 : romData <= 32'h61742065;
      11'b11101011011 : romData <= 32'h74656772;
      11'b11101011100 : romData <= 32'h74656220;
      11'b11101011101 : romData <= 32'h6E656577;
      11'b11101011110 : romData <= 32'h52445320;
      11'b11101011111 : romData <= 32'h28206D61;
      11'b11101100000 : romData <= 32'h61666564;
      11'b11101100001 : romData <= 32'h29746C75;
      11'b11101100010 : romData <= 32'h646E6120;
      11'b11101100011 : romData <= 32'h616C4620;
      11'b11101100100 : romData <= 32'h000A6873;
      11'b11101100101 : romData <= 32'h50206D2A;
      11'b11101100110 : romData <= 32'h6F667265;
      11'b11101100111 : romData <= 32'h73206D72;
      11'b11101101000 : romData <= 32'h6C706D69;
      11'b11101101001 : romData <= 32'h44532065;
      11'b11101101010 : romData <= 32'h206D6152;
      11'b11101101011 : romData <= 32'h636D656D;
      11'b11101101100 : romData <= 32'h6B636568;
      11'b11101101101 : romData <= 32'h732A000A;
      11'b11101101110 : romData <= 32'h65684320;
      11'b11101101111 : romData <= 32'h53206B63;
      11'b11101110000 : romData <= 32'h662D4950;
      11'b11101110001 : romData <= 32'h6873616C;
      11'b11101110010 : romData <= 32'h69686320;
      11'b11101110011 : romData <= 32'h2A000A70;
      11'b11101110100 : romData <= 32'h72452065;
      11'b11101110101 : romData <= 32'h20657361;
      11'b11101110110 : romData <= 32'h2D495053;
      11'b11101110111 : romData <= 32'h73616C66;
      11'b11101111000 : romData <= 32'h68632068;
      11'b11101111001 : romData <= 32'h000A7069;
      11'b11101111010 : romData <= 32'h5220722A;
      11'b11101111011 : romData <= 32'h70206E75;
      11'b11101111100 : romData <= 32'h72676F72;
      11'b11101111101 : romData <= 32'h69206D61;
      11'b11101111110 : romData <= 32'h5053206E;
      11'b11101111111 : romData <= 32'h6C662D49;
      11'b11110000000 : romData <= 32'h0A687361;
      11'b11110000001 : romData <= 32'h20662A00;
      11'b11110000010 : romData <= 32'h726F7453;
      11'b11110000011 : romData <= 32'h72702065;
      11'b11110000100 : romData <= 32'h6172676F;
      11'b11110000101 : romData <= 32'h6F6C206D;
      11'b11110000110 : romData <= 32'h64656461;
      11'b11110000111 : romData <= 32'h206E6920;
      11'b11110001000 : romData <= 32'h41524453;
      11'b11110001001 : romData <= 32'h6F74204D;
      11'b11110001010 : romData <= 32'h49505320;
      11'b11110001011 : romData <= 32'h616C462D;
      11'b11110001100 : romData <= 32'h000A6873;
      11'b11110001101 : romData <= 32'h4320632A;
      11'b11110001110 : romData <= 32'h61706D6F;
      11'b11110001111 : romData <= 32'h70206572;
      11'b11110010000 : romData <= 32'h72676F72;
      11'b11110010001 : romData <= 32'h6C206D61;
      11'b11110010010 : romData <= 32'h6564616F;
      11'b11110010011 : romData <= 32'h6E692064;
      11'b11110010100 : romData <= 32'h52445320;
      11'b11110010101 : romData <= 32'h77204D41;
      11'b11110010110 : romData <= 32'h20687469;
      11'b11110010111 : romData <= 32'h2D495053;
      11'b11110011000 : romData <= 32'h73616C46;
      11'b11110011001 : romData <= 32'h2A000A68;
      11'b11110011010 : romData <= 32'h68542068;
      11'b11110011011 : romData <= 32'h68207369;
      11'b11110011100 : romData <= 32'h73706C65;
      11'b11110011101 : romData <= 32'h65657263;
      11'b11110011110 : romData <= 32'h000A0A6E;
      11'b11110011111 : romData <= 32'hEFBEADDE;
      11'b11110100000 : romData <= 32'h01000000;
      11'b11110100001 : romData <= 32'h02000000;
      11'b11110100010 : romData <= 32'h03000000;
      11'b11110100011 : romData <= 32'h04000000;
      11'b11110100100 : romData <= 32'h05000000;
      11'b11110100101 : romData <= 32'h06000000;
      11'b11110100110 : romData <= 32'h07000000;
      11'b11110100111 : romData <= 32'hC21C00F0;
      11'b11110101000 : romData <= 32'hD91C00F0;
      11'b11110101001 : romData <= 32'h001D00F0;
      11'b11110101010 : romData <= 32'h231D00F0;
      11'b11110101011 : romData <= 32'h3D1D00F0;
      11'b11110101100 : romData <= 32'h601D00F0;
      11'b11110101101 : romData <= 32'h941D00F0;
      11'b11110101110 : romData <= 32'hB61D00F0;
      11'b11110101111 : romData <= 32'hCF1D00F0;
      11'b11110110000 : romData <= 32'hE81D00F0;
      11'b11110110001 : romData <= 32'h051E00F0;
      11'b11110110010 : romData <= 32'h341E00F0;
      11'b11110110011 : romData <= 32'h671E00F0;
      11'b11110110101 : romData <= 32'h10000000;
      11'b11110110111 : romData <= 32'h00527A01;
      11'b11110111000 : romData <= 32'h01097C04;
      11'b11110111001 : romData <= 32'h00010D1B;
      11'b11110111010 : romData <= 32'h14000000;
      11'b11110111011 : romData <= 32'h18000000;
      11'b11110111100 : romData <= 32'hBCF8FFFF;
      11'b11110111101 : romData <= 32'h14000000;
      11'b11110111110 : romData <= 32'h09094100;
      11'b11110111111 : romData <= 32'h0000000D;
      default : romData <= 32'd0;
    endcase

endmodule

